`timescale 1ns/1ps

module vga(clk);
   input clk;
   wire [16-1:0] result[1024-1:0];
   reg [144-1:0] memory [1024-1:0];
   reg [32-1:0]  counter;
   wire 	 vb [1024-1:0];
   reg [16-1:0]  graphicsMem [1024-1:0];

   integer 	 write_file;
   integer 	 read_data;
   
   generator gn817 (memory[817], 817, counter, result[817], vb[817]);
   generator gn620 (memory[620], 620, counter, result[620], vb[620]);
   generator gn293 (memory[293], 293, counter, result[293], vb[293]);
   generator gn712 (memory[712], 712, counter, result[712], vb[712]);
   generator gn35 (memory[35], 35, counter, result[35], vb[35]);
   generator gn673 (memory[673], 673, counter, result[673], vb[673]);
   generator gn601 (memory[601], 601, counter, result[601], vb[601]);
   generator gn517 (memory[517], 517, counter, result[517], vb[517]);
   generator gn200 (memory[200], 200, counter, result[200], vb[200]);
   generator gn431 (memory[431], 431, counter, result[431], vb[431]);
   generator gn950 (memory[950], 950, counter, result[950], vb[950]);
   generator gn183 (memory[183], 183, counter, result[183], vb[183]);
   generator gn276 (memory[276], 276, counter, result[276], vb[276]);
   generator gn441 (memory[441], 441, counter, result[441], vb[441]);
   generator gn584 (memory[584], 584, counter, result[584], vb[584]);
   generator gn467 (memory[467], 467, counter, result[467], vb[467]);
   generator gn839 (memory[839], 839, counter, result[839], vb[839]);
   generator gn104 (memory[104], 104, counter, result[104], vb[104]);
   generator gn331 (memory[331], 331, counter, result[331], vb[331]);
   generator gn529 (memory[529], 529, counter, result[529], vb[529]);
   generator gn49 (memory[49], 49, counter, result[49], vb[49]);
   generator gn22 (memory[22], 22, counter, result[22], vb[22]);
   generator gn451 (memory[451], 451, counter, result[451], vb[451]);
   generator gn1008 (memory[1008], 1008, counter, result[1008], vb[1008]);
   generator gn685 (memory[685], 685, counter, result[685], vb[685]);
   generator gn297 (memory[297], 297, counter, result[297], vb[297]);
   generator gn343 (memory[343], 343, counter, result[343], vb[343]);
   generator gn579 (memory[579], 579, counter, result[579], vb[579]);
   generator gn701 (memory[701], 701, counter, result[701], vb[701]);
   generator gn1012 (memory[1012], 1012, counter, result[1012], vb[1012]);
   generator gn1013 (memory[1013], 1013, counter, result[1013], vb[1013]);
   generator gn439 (memory[439], 439, counter, result[439], vb[439]);
   generator gn391 (memory[391], 391, counter, result[391], vb[391]);
   generator gn981 (memory[981], 981, counter, result[981], vb[981]);
   generator gn889 (memory[889], 889, counter, result[889], vb[889]);
   generator gn305 (memory[305], 305, counter, result[305], vb[305]);
   generator gn105 (memory[105], 105, counter, result[105], vb[105]);
   generator gn187 (memory[187], 187, counter, result[187], vb[187]);
   generator gn616 (memory[616], 616, counter, result[616], vb[616]);
   generator gn569 (memory[569], 569, counter, result[569], vb[569]);
   generator gn154 (memory[154], 154, counter, result[154], vb[154]);
   generator gn476 (memory[476], 476, counter, result[476], vb[476]);
   generator gn54 (memory[54], 54, counter, result[54], vb[54]);
   generator gn468 (memory[468], 468, counter, result[468], vb[468]);
   generator gn629 (memory[629], 629, counter, result[629], vb[629]);
   generator gn648 (memory[648], 648, counter, result[648], vb[648]);
   generator gn100 (memory[100], 100, counter, result[100], vb[100]);
   generator gn850 (memory[850], 850, counter, result[850], vb[850]);
   generator gn888 (memory[888], 888, counter, result[888], vb[888]);
   generator gn376 (memory[376], 376, counter, result[376], vb[376]);
   generator gn434 (memory[434], 434, counter, result[434], vb[434]);
   generator gn955 (memory[955], 955, counter, result[955], vb[955]);
   generator gn273 (memory[273], 273, counter, result[273], vb[273]);
   generator gn463 (memory[463], 463, counter, result[463], vb[463]);
   generator gn157 (memory[157], 157, counter, result[157], vb[157]);
   generator gn635 (memory[635], 635, counter, result[635], vb[635]);
   generator gn968 (memory[968], 968, counter, result[968], vb[968]);
   generator gn291 (memory[291], 291, counter, result[291], vb[291]);
   generator gn493 (memory[493], 493, counter, result[493], vb[493]);
   generator gn934 (memory[934], 934, counter, result[934], vb[934]);
   generator gn113 (memory[113], 113, counter, result[113], vb[113]);
   generator gn289 (memory[289], 289, counter, result[289], vb[289]);
   generator gn651 (memory[651], 651, counter, result[651], vb[651]);
   generator gn38 (memory[38], 38, counter, result[38], vb[38]);
   generator gn900 (memory[900], 900, counter, result[900], vb[900]);
   generator gn724 (memory[724], 724, counter, result[724], vb[724]);
   generator gn292 (memory[292], 292, counter, result[292], vb[292]);
   generator gn713 (memory[713], 713, counter, result[713], vb[713]);
   generator gn162 (memory[162], 162, counter, result[162], vb[162]);
   generator gn102 (memory[102], 102, counter, result[102], vb[102]);
   generator gn248 (memory[248], 248, counter, result[248], vb[248]);
   generator gn284 (memory[284], 284, counter, result[284], vb[284]);
   generator gn76 (memory[76], 76, counter, result[76], vb[76]);
   generator gn811 (memory[811], 811, counter, result[811], vb[811]);
   generator gn473 (memory[473], 473, counter, result[473], vb[473]);
   generator gn645 (memory[645], 645, counter, result[645], vb[645]);
   generator gn678 (memory[678], 678, counter, result[678], vb[678]);
   generator gn650 (memory[650], 650, counter, result[650], vb[650]);
   generator gn985 (memory[985], 985, counter, result[985], vb[985]);
   generator gn769 (memory[769], 769, counter, result[769], vb[769]);
   generator gn536 (memory[536], 536, counter, result[536], vb[536]);
   generator gn935 (memory[935], 935, counter, result[935], vb[935]);
   generator gn406 (memory[406], 406, counter, result[406], vb[406]);
   generator gn423 (memory[423], 423, counter, result[423], vb[423]);
   generator gn1021 (memory[1021], 1021, counter, result[1021], vb[1021]);
   generator gn967 (memory[967], 967, counter, result[967], vb[967]);
   generator gn37 (memory[37], 37, counter, result[37], vb[37]);
   generator gn1023 (memory[1023], 1023, counter, result[1023], vb[1023]);
   generator gn840 (memory[840], 840, counter, result[840], vb[840]);
   generator gn345 (memory[345], 345, counter, result[345], vb[345]);
   generator gn774 (memory[774], 774, counter, result[774], vb[774]);
   generator gn45 (memory[45], 45, counter, result[45], vb[45]);
   generator gn181 (memory[181], 181, counter, result[181], vb[181]);
   generator gn412 (memory[412], 412, counter, result[412], vb[412]);
   generator gn554 (memory[554], 554, counter, result[554], vb[554]);
   generator gn311 (memory[311], 311, counter, result[311], vb[311]);
   generator gn384 (memory[384], 384, counter, result[384], vb[384]);
   generator gn137 (memory[137], 137, counter, result[137], vb[137]);
   generator gn956 (memory[956], 956, counter, result[956], vb[956]);
   generator gn808 (memory[808], 808, counter, result[808], vb[808]);
   generator gn469 (memory[469], 469, counter, result[469], vb[469]);
   generator gn46 (memory[46], 46, counter, result[46], vb[46]);
   generator gn542 (memory[542], 542, counter, result[542], vb[542]);
   generator gn675 (memory[675], 675, counter, result[675], vb[675]);
   generator gn775 (memory[775], 775, counter, result[775], vb[775]);
   generator gn921 (memory[921], 921, counter, result[921], vb[921]);
   generator gn156 (memory[156], 156, counter, result[156], vb[156]);
   generator gn462 (memory[462], 462, counter, result[462], vb[462]);
   generator gn903 (memory[903], 903, counter, result[903], vb[903]);
   generator gn127 (memory[127], 127, counter, result[127], vb[127]);
   generator gn454 (memory[454], 454, counter, result[454], vb[454]);
   generator gn730 (memory[730], 730, counter, result[730], vb[730]);
   generator gn40 (memory[40], 40, counter, result[40], vb[40]);
   generator gn595 (memory[595], 595, counter, result[595], vb[595]);
   generator gn931 (memory[931], 931, counter, result[931], vb[931]);
   generator gn617 (memory[617], 617, counter, result[617], vb[617]);
   generator gn298 (memory[298], 298, counter, result[298], vb[298]);
   generator gn2 (memory[2], 2, counter, result[2], vb[2]);
   generator gn315 (memory[315], 315, counter, result[315], vb[315]);
   generator gn942 (memory[942], 942, counter, result[942], vb[942]);
   generator gn394 (memory[394], 394, counter, result[394], vb[394]);
   generator gn729 (memory[729], 729, counter, result[729], vb[729]);
   generator gn503 (memory[503], 503, counter, result[503], vb[503]);
   generator gn122 (memory[122], 122, counter, result[122], vb[122]);
   generator gn97 (memory[97], 97, counter, result[97], vb[97]);
   generator gn225 (memory[225], 225, counter, result[225], vb[225]);
   generator gn470 (memory[470], 470, counter, result[470], vb[470]);
   generator gn717 (memory[717], 717, counter, result[717], vb[717]);
   generator gn84 (memory[84], 84, counter, result[84], vb[84]);
   generator gn109 (memory[109], 109, counter, result[109], vb[109]);
   generator gn649 (memory[649], 649, counter, result[649], vb[649]);
   generator gn797 (memory[797], 797, counter, result[797], vb[797]);
   generator gn692 (memory[692], 692, counter, result[692], vb[692]);
   generator gn1005 (memory[1005], 1005, counter, result[1005], vb[1005]);
   generator gn247 (memory[247], 247, counter, result[247], vb[247]);
   generator gn844 (memory[844], 844, counter, result[844], vb[844]);
   generator gn933 (memory[933], 933, counter, result[933], vb[933]);
   generator gn31 (memory[31], 31, counter, result[31], vb[31]);
   generator gn705 (memory[705], 705, counter, result[705], vb[705]);
   generator gn904 (memory[904], 904, counter, result[904], vb[904]);
   generator gn1 (memory[1], 1, counter, result[1], vb[1]);
   generator gn101 (memory[101], 101, counter, result[101], vb[101]);
   generator gn23 (memory[23], 23, counter, result[23], vb[23]);
   generator gn515 (memory[515], 515, counter, result[515], vb[515]);
   generator gn943 (memory[943], 943, counter, result[943], vb[943]);
   generator gn27 (memory[27], 27, counter, result[27], vb[27]);
   generator gn758 (memory[758], 758, counter, result[758], vb[758]);
   generator gn203 (memory[203], 203, counter, result[203], vb[203]);
   generator gn372 (memory[372], 372, counter, result[372], vb[372]);
   generator gn992 (memory[992], 992, counter, result[992], vb[992]);
   generator gn175 (memory[175], 175, counter, result[175], vb[175]);
   generator gn498 (memory[498], 498, counter, result[498], vb[498]);
   generator gn519 (memory[519], 519, counter, result[519], vb[519]);
   generator gn228 (memory[228], 228, counter, result[228], vb[228]);
   generator gn874 (memory[874], 874, counter, result[874], vb[874]);
   generator gn897 (memory[897], 897, counter, result[897], vb[897]);
   generator gn777 (memory[777], 777, counter, result[777], vb[777]);
   generator gn731 (memory[731], 731, counter, result[731], vb[731]);
   generator gn513 (memory[513], 513, counter, result[513], vb[513]);
   generator gn668 (memory[668], 668, counter, result[668], vb[668]);
   generator gn546 (memory[546], 546, counter, result[546], vb[546]);
   generator gn671 (memory[671], 671, counter, result[671], vb[671]);
   generator gn1018 (memory[1018], 1018, counter, result[1018], vb[1018]);
   generator gn226 (memory[226], 226, counter, result[226], vb[226]);
   generator gn218 (memory[218], 218, counter, result[218], vb[218]);
   generator gn9 (memory[9], 9, counter, result[9], vb[9]);
   generator gn405 (memory[405], 405, counter, result[405], vb[405]);
   generator gn737 (memory[737], 737, counter, result[737], vb[737]);
   generator gn359 (memory[359], 359, counter, result[359], vb[359]);
   generator gn908 (memory[908], 908, counter, result[908], vb[908]);
   generator gn804 (memory[804], 804, counter, result[804], vb[804]);
   generator gn161 (memory[161], 161, counter, result[161], vb[161]);
   generator gn784 (memory[784], 784, counter, result[784], vb[784]);
   generator gn208 (memory[208], 208, counter, result[208], vb[208]);
   generator gn929 (memory[929], 929, counter, result[929], vb[929]);
   generator gn680 (memory[680], 680, counter, result[680], vb[680]);
   generator gn504 (memory[504], 504, counter, result[504], vb[504]);
   generator gn590 (memory[590], 590, counter, result[590], vb[590]);
   generator gn361 (memory[361], 361, counter, result[361], vb[361]);
   generator gn899 (memory[899], 899, counter, result[899], vb[899]);
   generator gn711 (memory[711], 711, counter, result[711], vb[711]);
   generator gn374 (memory[374], 374, counter, result[374], vb[374]);
   generator gn354 (memory[354], 354, counter, result[354], vb[354]);
   generator gn172 (memory[172], 172, counter, result[172], vb[172]);
   generator gn789 (memory[789], 789, counter, result[789], vb[789]);
   generator gn344 (memory[344], 344, counter, result[344], vb[344]);
   generator gn255 (memory[255], 255, counter, result[255], vb[255]);
   generator gn336 (memory[336], 336, counter, result[336], vb[336]);
   generator gn571 (memory[571], 571, counter, result[571], vb[571]);
   generator gn858 (memory[858], 858, counter, result[858], vb[858]);
   generator gn316 (memory[316], 316, counter, result[316], vb[316]);
   generator gn232 (memory[232], 232, counter, result[232], vb[232]);
   generator gn767 (memory[767], 767, counter, result[767], vb[767]);
   generator gn220 (memory[220], 220, counter, result[220], vb[220]);
   generator gn939 (memory[939], 939, counter, result[939], vb[939]);
   generator gn977 (memory[977], 977, counter, result[977], vb[977]);
   generator gn174 (memory[174], 174, counter, result[174], vb[174]);
   generator gn360 (memory[360], 360, counter, result[360], vb[360]);
   generator gn303 (memory[303], 303, counter, result[303], vb[303]);
   generator gn998 (memory[998], 998, counter, result[998], vb[998]);
   generator gn93 (memory[93], 93, counter, result[93], vb[93]);
   generator gn204 (memory[204], 204, counter, result[204], vb[204]);
   generator gn90 (memory[90], 90, counter, result[90], vb[90]);
   generator gn854 (memory[854], 854, counter, result[854], vb[854]);
   generator gn395 (memory[395], 395, counter, result[395], vb[395]);
   generator gn237 (memory[237], 237, counter, result[237], vb[237]);
   generator gn823 (memory[823], 823, counter, result[823], vb[823]);
   generator gn263 (memory[263], 263, counter, result[263], vb[263]);
   generator gn990 (memory[990], 990, counter, result[990], vb[990]);
   generator gn560 (memory[560], 560, counter, result[560], vb[560]);
   generator gn734 (memory[734], 734, counter, result[734], vb[734]);
   generator gn852 (memory[852], 852, counter, result[852], vb[852]);
   generator gn885 (memory[885], 885, counter, result[885], vb[885]);
   generator gn790 (memory[790], 790, counter, result[790], vb[790]);
   generator gn318 (memory[318], 318, counter, result[318], vb[318]);
   generator gn941 (memory[941], 941, counter, result[941], vb[941]);
   generator gn766 (memory[766], 766, counter, result[766], vb[766]);
   generator gn791 (memory[791], 791, counter, result[791], vb[791]);
   generator gn526 (memory[526], 526, counter, result[526], vb[526]);
   generator gn953 (memory[953], 953, counter, result[953], vb[953]);
   generator gn991 (memory[991], 991, counter, result[991], vb[991]);
   generator gn785 (memory[785], 785, counter, result[785], vb[785]);
   generator gn902 (memory[902], 902, counter, result[902], vb[902]);
   generator gn975 (memory[975], 975, counter, result[975], vb[975]);
   generator gn857 (memory[857], 857, counter, result[857], vb[857]);
   generator gn15 (memory[15], 15, counter, result[15], vb[15]);
   generator gn495 (memory[495], 495, counter, result[495], vb[495]);
   generator gn160 (memory[160], 160, counter, result[160], vb[160]);
   generator gn346 (memory[346], 346, counter, result[346], vb[346]);
   generator gn786 (memory[786], 786, counter, result[786], vb[786]);
   generator gn656 (memory[656], 656, counter, result[656], vb[656]);
   generator gn29 (memory[29], 29, counter, result[29], vb[29]);
   generator gn142 (memory[142], 142, counter, result[142], vb[142]);
   generator gn756 (memory[756], 756, counter, result[756], vb[756]);
   generator gn572 (memory[572], 572, counter, result[572], vb[572]);
   generator gn793 (memory[793], 793, counter, result[793], vb[793]);
   generator gn715 (memory[715], 715, counter, result[715], vb[715]);
   generator gn838 (memory[838], 838, counter, result[838], vb[838]);
   generator gn1010 (memory[1010], 1010, counter, result[1010], vb[1010]);
   generator gn832 (memory[832], 832, counter, result[832], vb[832]);
   generator gn433 (memory[433], 433, counter, result[433], vb[433]);
   generator gn720 (memory[720], 720, counter, result[720], vb[720]);
   generator gn851 (memory[851], 851, counter, result[851], vb[851]);
   generator gn566 (memory[566], 566, counter, result[566], vb[566]);
   generator gn849 (memory[849], 849, counter, result[849], vb[849]);
   generator gn231 (memory[231], 231, counter, result[231], vb[231]);
   generator gn216 (memory[216], 216, counter, result[216], vb[216]);
   generator gn794 (memory[794], 794, counter, result[794], vb[794]);
   generator gn474 (memory[474], 474, counter, result[474], vb[474]);
   generator gn841 (memory[841], 841, counter, result[841], vb[841]);
   generator gn171 (memory[171], 171, counter, result[171], vb[171]);
   generator gn927 (memory[927], 927, counter, result[927], vb[927]);
   generator gn690 (memory[690], 690, counter, result[690], vb[690]);
   generator gn835 (memory[835], 835, counter, result[835], vb[835]);
   generator gn383 (memory[383], 383, counter, result[383], vb[383]);
   generator gn99 (memory[99], 99, counter, result[99], vb[99]);
   generator gn613 (memory[613], 613, counter, result[613], vb[613]);
   generator gn0 (memory[0], 0, counter, result[0], vb[0]);
   generator gn780 (memory[780], 780, counter, result[780], vb[780]);
   generator gn482 (memory[482], 482, counter, result[482], vb[482]);
   generator gn347 (memory[347], 347, counter, result[347], vb[347]);
   generator gn337 (memory[337], 337, counter, result[337], vb[337]);
   generator gn938 (memory[938], 938, counter, result[938], vb[938]);
   generator gn700 (memory[700], 700, counter, result[700], vb[700]);
   generator gn615 (memory[615], 615, counter, result[615], vb[615]);
   generator gn487 (memory[487], 487, counter, result[487], vb[487]);
   generator gn159 (memory[159], 159, counter, result[159], vb[159]);
   generator gn322 (memory[322], 322, counter, result[322], vb[322]);
   generator gn96 (memory[96], 96, counter, result[96], vb[96]);
   generator gn708 (memory[708], 708, counter, result[708], vb[708]);
   generator gn703 (memory[703], 703, counter, result[703], vb[703]);
   generator gn271 (memory[271], 271, counter, result[271], vb[271]);
   generator gn867 (memory[867], 867, counter, result[867], vb[867]);
   generator gn274 (memory[274], 274, counter, result[274], vb[274]);
   generator gn637 (memory[637], 637, counter, result[637], vb[637]);
   generator gn98 (memory[98], 98, counter, result[98], vb[98]);
   generator gn327 (memory[327], 327, counter, result[327], vb[327]);
   generator gn864 (memory[864], 864, counter, result[864], vb[864]);
   generator gn779 (memory[779], 779, counter, result[779], vb[779]);
   generator gn1020 (memory[1020], 1020, counter, result[1020], vb[1020]);
   generator gn866 (memory[866], 866, counter, result[866], vb[866]);
   generator gn414 (memory[414], 414, counter, result[414], vb[414]);
   generator gn432 (memory[432], 432, counter, result[432], vb[432]);
   generator gn805 (memory[805], 805, counter, result[805], vb[805]);
   generator gn833 (memory[833], 833, counter, result[833], vb[833]);
   generator gn143 (memory[143], 143, counter, result[143], vb[143]);
   generator gn633 (memory[633], 633, counter, result[633], vb[633]);
   generator gn847 (memory[847], 847, counter, result[847], vb[847]);
   generator gn449 (memory[449], 449, counter, result[449], vb[449]);
   generator gn746 (memory[746], 746, counter, result[746], vb[746]);
   generator gn81 (memory[81], 81, counter, result[81], vb[81]);
   generator gn642 (memory[642], 642, counter, result[642], vb[642]);
   generator gn599 (memory[599], 599, counter, result[599], vb[599]);
   generator gn920 (memory[920], 920, counter, result[920], vb[920]);
   generator gn267 (memory[267], 267, counter, result[267], vb[267]);
   generator gn557 (memory[557], 557, counter, result[557], vb[557]);
   generator gn951 (memory[951], 951, counter, result[951], vb[951]);
   generator gn883 (memory[883], 883, counter, result[883], vb[883]);
   generator gn585 (memory[585], 585, counter, result[585], vb[585]);
   generator gn120 (memory[120], 120, counter, result[120], vb[120]);
   generator gn188 (memory[188], 188, counter, result[188], vb[188]);
   generator gn3 (memory[3], 3, counter, result[3], vb[3]);
   generator gn600 (memory[600], 600, counter, result[600], vb[600]);
   generator gn676 (memory[676], 676, counter, result[676], vb[676]);
   generator gn916 (memory[916], 916, counter, result[916], vb[916]);
   generator gn444 (memory[444], 444, counter, result[444], vb[444]);
   generator gn80 (memory[80], 80, counter, result[80], vb[80]);
   generator gn223 (memory[223], 223, counter, result[223], vb[223]);
   generator gn568 (memory[568], 568, counter, result[568], vb[568]);
   generator gn295 (memory[295], 295, counter, result[295], vb[295]);
   generator gn438 (memory[438], 438, counter, result[438], vb[438]);
   generator gn402 (memory[402], 402, counter, result[402], vb[402]);
   generator gn755 (memory[755], 755, counter, result[755], vb[755]);
   generator gn26 (memory[26], 26, counter, result[26], vb[26]);
   generator gn69 (memory[69], 69, counter, result[69], vb[69]);
   generator gn550 (memory[550], 550, counter, result[550], vb[550]);
   generator gn828 (memory[828], 828, counter, result[828], vb[828]);
   generator gn329 (memory[329], 329, counter, result[329], vb[329]);
   generator gn340 (memory[340], 340, counter, result[340], vb[340]);
   generator gn198 (memory[198], 198, counter, result[198], vb[198]);
   generator gn625 (memory[625], 625, counter, result[625], vb[625]);
   generator gn268 (memory[268], 268, counter, result[268], vb[268]);
   generator gn68 (memory[68], 68, counter, result[68], vb[68]);
   generator gn456 (memory[456], 456, counter, result[456], vb[456]);
   generator gn338 (memory[338], 338, counter, result[338], vb[338]);
   generator gn310 (memory[310], 310, counter, result[310], vb[310]);
   generator gn499 (memory[499], 499, counter, result[499], vb[499]);
   generator gn508 (memory[508], 508, counter, result[508], vb[508]);
   generator gn13 (memory[13], 13, counter, result[13], vb[13]);
   generator gn108 (memory[108], 108, counter, result[108], vb[108]);
   generator gn400 (memory[400], 400, counter, result[400], vb[400]);
   generator gn34 (memory[34], 34, counter, result[34], vb[34]);
   generator gn119 (memory[119], 119, counter, result[119], vb[119]);
   generator gn646 (memory[646], 646, counter, result[646], vb[646]);
   generator gn528 (memory[528], 528, counter, result[528], vb[528]);
   generator gn328 (memory[328], 328, counter, result[328], vb[328]);
   generator gn604 (memory[604], 604, counter, result[604], vb[604]);
   generator gn124 (memory[124], 124, counter, result[124], vb[124]);
   generator gn527 (memory[527], 527, counter, result[527], vb[527]);
   generator gn472 (memory[472], 472, counter, result[472], vb[472]);
   generator gn207 (memory[207], 207, counter, result[207], vb[207]);
   generator gn75 (memory[75], 75, counter, result[75], vb[75]);
   generator gn699 (memory[699], 699, counter, result[699], vb[699]);
   generator gn241 (memory[241], 241, counter, result[241], vb[241]);
   generator gn578 (memory[578], 578, counter, result[578], vb[578]);
   generator gn73 (memory[73], 73, counter, result[73], vb[73]);
   generator gn996 (memory[996], 996, counter, result[996], vb[996]);
   generator gn130 (memory[130], 130, counter, result[130], vb[130]);
   generator gn121 (memory[121], 121, counter, result[121], vb[121]);
   generator gn984 (memory[984], 984, counter, result[984], vb[984]);
   generator gn86 (memory[86], 86, counter, result[86], vb[86]);
   generator gn63 (memory[63], 63, counter, result[63], vb[63]);
   generator gn597 (memory[597], 597, counter, result[597], vb[597]);
   generator gn684 (memory[684], 684, counter, result[684], vb[684]);
   generator gn184 (memory[184], 184, counter, result[184], vb[184]);
   generator gn14 (memory[14], 14, counter, result[14], vb[14]);
   generator gn326 (memory[326], 326, counter, result[326], vb[326]);
   generator gn365 (memory[365], 365, counter, result[365], vb[365]);
   generator gn845 (memory[845], 845, counter, result[845], vb[845]);
   generator gn380 (memory[380], 380, counter, result[380], vb[380]);
   generator gn370 (memory[370], 370, counter, result[370], vb[370]);
   generator gn25 (memory[25], 25, counter, result[25], vb[25]);
   generator gn562 (memory[562], 562, counter, result[562], vb[562]);
   generator gn364 (memory[364], 364, counter, result[364], vb[364]);
   generator gn919 (memory[919], 919, counter, result[919], vb[919]);
   generator gn702 (memory[702], 702, counter, result[702], vb[702]);
   generator gn424 (memory[424], 424, counter, result[424], vb[424]);
   generator gn362 (memory[362], 362, counter, result[362], vb[362]);
   generator gn693 (memory[693], 693, counter, result[693], vb[693]);
   generator gn957 (memory[957], 957, counter, result[957], vb[957]);
   generator gn420 (memory[420], 420, counter, result[420], vb[420]);
   generator gn825 (memory[825], 825, counter, result[825], vb[825]);
   generator gn398 (memory[398], 398, counter, result[398], vb[398]);
   generator gn94 (memory[94], 94, counter, result[94], vb[94]);
   generator gn138 (memory[138], 138, counter, result[138], vb[138]);
   generator gn489 (memory[489], 489, counter, result[489], vb[489]);
   generator gn773 (memory[773], 773, counter, result[773], vb[773]);
   generator gn771 (memory[771], 771, counter, result[771], vb[771]);
   generator gn357 (memory[357], 357, counter, result[357], vb[357]);
   generator gn843 (memory[843], 843, counter, result[843], vb[843]);
   generator gn707 (memory[707], 707, counter, result[707], vb[707]);
   generator gn483 (memory[483], 483, counter, result[483], vb[483]);
   generator gn638 (memory[638], 638, counter, result[638], vb[638]);
   generator gn182 (memory[182], 182, counter, result[182], vb[182]);
   generator gn43 (memory[43], 43, counter, result[43], vb[43]);
   generator gn619 (memory[619], 619, counter, result[619], vb[619]);
   generator gn275 (memory[275], 275, counter, result[275], vb[275]);
   generator gn453 (memory[453], 453, counter, result[453], vb[453]);
   generator gn719 (memory[719], 719, counter, result[719], vb[719]);
   generator gn577 (memory[577], 577, counter, result[577], vb[577]);
   generator gn588 (memory[588], 588, counter, result[588], vb[588]);
   generator gn926 (memory[926], 926, counter, result[926], vb[926]);
   generator gn622 (memory[622], 622, counter, result[622], vb[622]);
   generator gn309 (memory[309], 309, counter, result[309], vb[309]);
   generator gn873 (memory[873], 873, counter, result[873], vb[873]);
   generator gn1004 (memory[1004], 1004, counter, result[1004], vb[1004]);
   generator gn681 (memory[681], 681, counter, result[681], vb[681]);
   generator gn792 (memory[792], 792, counter, result[792], vb[792]);
   generator gn56 (memory[56], 56, counter, result[56], vb[56]);
   generator gn537 (memory[537], 537, counter, result[537], vb[537]);
   generator gn466 (memory[466], 466, counter, result[466], vb[466]);
   generator gn547 (memory[547], 547, counter, result[547], vb[547]);
   generator gn575 (memory[575], 575, counter, result[575], vb[575]);
   generator gn661 (memory[661], 661, counter, result[661], vb[661]);
   generator gn753 (memory[753], 753, counter, result[753], vb[753]);
   generator gn33 (memory[33], 33, counter, result[33], vb[33]);
   generator gn603 (memory[603], 603, counter, result[603], vb[603]);
   generator gn728 (memory[728], 728, counter, result[728], vb[728]);
   generator gn683 (memory[683], 683, counter, result[683], vb[683]);
   generator gn66 (memory[66], 66, counter, result[66], vb[66]);
   generator gn135 (memory[135], 135, counter, result[135], vb[135]);
   generator gn219 (memory[219], 219, counter, result[219], vb[219]);
   generator gn229 (memory[229], 229, counter, result[229], vb[229]);
   generator gn389 (memory[389], 389, counter, result[389], vb[389]);
   generator gn725 (memory[725], 725, counter, result[725], vb[725]);
   generator gn260 (memory[260], 260, counter, result[260], vb[260]);
   generator gn923 (memory[923], 923, counter, result[923], vb[923]);
   generator gn189 (memory[189], 189, counter, result[189], vb[189]);
   generator gn733 (memory[733], 733, counter, result[733], vb[733]);
   generator gn227 (memory[227], 227, counter, result[227], vb[227]);
   generator gn659 (memory[659], 659, counter, result[659], vb[659]);
   generator gn787 (memory[787], 787, counter, result[787], vb[787]);
   generator gn679 (memory[679], 679, counter, result[679], vb[679]);
   generator gn492 (memory[492], 492, counter, result[492], vb[492]);
   generator gn732 (memory[732], 732, counter, result[732], vb[732]);
   generator gn279 (memory[279], 279, counter, result[279], vb[279]);
   generator gn893 (memory[893], 893, counter, result[893], vb[893]);
   generator gn802 (memory[802], 802, counter, result[802], vb[802]);
   generator gn30 (memory[30], 30, counter, result[30], vb[30]);
   generator gn1000 (memory[1000], 1000, counter, result[1000], vb[1000]);
   generator gn949 (memory[949], 949, counter, result[949], vb[949]);
   generator gn570 (memory[570], 570, counter, result[570], vb[570]);
   generator gn634 (memory[634], 634, counter, result[634], vb[634]);
   generator gn464 (memory[464], 464, counter, result[464], vb[464]);
   generator gn144 (memory[144], 144, counter, result[144], vb[144]);
   generator gn522 (memory[522], 522, counter, result[522], vb[522]);
   generator gn1014 (memory[1014], 1014, counter, result[1014], vb[1014]);
   generator gn11 (memory[11], 11, counter, result[11], vb[11]);
   generator gn763 (memory[763], 763, counter, result[763], vb[763]);
   generator gn759 (memory[759], 759, counter, result[759], vb[759]);
   generator gn418 (memory[418], 418, counter, result[418], vb[418]);
   generator gn909 (memory[909], 909, counter, result[909], vb[909]);
   generator gn335 (memory[335], 335, counter, result[335], vb[335]);
   generator gn895 (memory[895], 895, counter, result[895], vb[895]);
   generator gn50 (memory[50], 50, counter, result[50], vb[50]);
   generator gn842 (memory[842], 842, counter, result[842], vb[842]);
   generator gn249 (memory[249], 249, counter, result[249], vb[249]);
   generator gn624 (memory[624], 624, counter, result[624], vb[624]);
   generator gn962 (memory[962], 962, counter, result[962], vb[962]);
   generator gn995 (memory[995], 995, counter, result[995], vb[995]);
   generator gn1019 (memory[1019], 1019, counter, result[1019], vb[1019]);
   generator gn16 (memory[16], 16, counter, result[16], vb[16]);
   generator gn12 (memory[12], 12, counter, result[12], vb[12]);
   generator gn17 (memory[17], 17, counter, result[17], vb[17]);
   generator gn290 (memory[290], 290, counter, result[290], vb[290]);
   generator gn770 (memory[770], 770, counter, result[770], vb[770]);
   generator gn299 (memory[299], 299, counter, result[299], vb[299]);
   generator gn698 (memory[698], 698, counter, result[698], vb[698]);
   generator gn913 (memory[913], 913, counter, result[913], vb[913]);
   generator gn153 (memory[153], 153, counter, result[153], vb[153]);
   generator gn349 (memory[349], 349, counter, result[349], vb[349]);
   generator gn521 (memory[521], 521, counter, result[521], vb[521]);
   generator gn605 (memory[605], 605, counter, result[605], vb[605]);
   generator gn915 (memory[915], 915, counter, result[915], vb[915]);
   generator gn59 (memory[59], 59, counter, result[59], vb[59]);
   generator gn627 (memory[627], 627, counter, result[627], vb[627]);
   generator gn125 (memory[125], 125, counter, result[125], vb[125]);
   generator gn381 (memory[381], 381, counter, result[381], vb[381]);
   generator gn74 (memory[74], 74, counter, result[74], vb[74]);
   generator gn691 (memory[691], 691, counter, result[691], vb[691]);
   generator gn917 (memory[917], 917, counter, result[917], vb[917]);
   generator gn288 (memory[288], 288, counter, result[288], vb[288]);
   generator gn740 (memory[740], 740, counter, result[740], vb[740]);
   generator gn325 (memory[325], 325, counter, result[325], vb[325]);
   generator gn567 (memory[567], 567, counter, result[567], vb[567]);
   generator gn1002 (memory[1002], 1002, counter, result[1002], vb[1002]);
   generator gn798 (memory[798], 798, counter, result[798], vb[798]);
   generator gn602 (memory[602], 602, counter, result[602], vb[602]);
   generator gn195 (memory[195], 195, counter, result[195], vb[195]);
   generator gn686 (memory[686], 686, counter, result[686], vb[686]);
   generator gn334 (memory[334], 334, counter, result[334], vb[334]);
   generator gn781 (memory[781], 781, counter, result[781], vb[781]);
   generator gn535 (memory[535], 535, counter, result[535], vb[535]);
   generator gn972 (memory[972], 972, counter, result[972], vb[972]);
   generator gn110 (memory[110], 110, counter, result[110], vb[110]);
   generator gn856 (memory[856], 856, counter, result[856], vb[856]);
   generator gn491 (memory[491], 491, counter, result[491], vb[491]);
   generator gn657 (memory[657], 657, counter, result[657], vb[657]);
   generator gn397 (memory[397], 397, counter, result[397], vb[397]);
   generator gn158 (memory[158], 158, counter, result[158], vb[158]);
   generator gn598 (memory[598], 598, counter, result[598], vb[598]);
   generator gn822 (memory[822], 822, counter, result[822], vb[822]);
   generator gn722 (memory[722], 722, counter, result[722], vb[722]);
   generator gn243 (memory[243], 243, counter, result[243], vb[243]);
   generator gn178 (memory[178], 178, counter, result[178], vb[178]);
   generator gn721 (memory[721], 721, counter, result[721], vb[721]);
   generator gn323 (memory[323], 323, counter, result[323], vb[323]);
   generator gn230 (memory[230], 230, counter, result[230], vb[230]);
   generator gn884 (memory[884], 884, counter, result[884], vb[884]);
   generator gn860 (memory[860], 860, counter, result[860], vb[860]);
   generator gn596 (memory[596], 596, counter, result[596], vb[596]);
   generator gn148 (memory[148], 148, counter, result[148], vb[148]);
   generator gn621 (memory[621], 621, counter, result[621], vb[621]);
   generator gn606 (memory[606], 606, counter, result[606], vb[606]);
   generator gn593 (memory[593], 593, counter, result[593], vb[593]);
   generator gn387 (memory[387], 387, counter, result[387], vb[387]);
   generator gn905 (memory[905], 905, counter, result[905], vb[905]);
   generator gn533 (memory[533], 533, counter, result[533], vb[533]);
   generator gn907 (memory[907], 907, counter, result[907], vb[907]);
   generator gn757 (memory[757], 757, counter, result[757], vb[757]);
   generator gn744 (memory[744], 744, counter, result[744], vb[744]);
   generator gn639 (memory[639], 639, counter, result[639], vb[639]);
   generator gn202 (memory[202], 202, counter, result[202], vb[202]);
   generator gn317 (memory[317], 317, counter, result[317], vb[317]);
   generator gn824 (memory[824], 824, counter, result[824], vb[824]);
   generator gn932 (memory[932], 932, counter, result[932], vb[932]);
   generator gn837 (memory[837], 837, counter, result[837], vb[837]);
   generator gn501 (memory[501], 501, counter, result[501], vb[501]);
   generator gn742 (memory[742], 742, counter, result[742], vb[742]);
   generator gn368 (memory[368], 368, counter, result[368], vb[368]);
   generator gn111 (memory[111], 111, counter, result[111], vb[111]);
   generator gn1001 (memory[1001], 1001, counter, result[1001], vb[1001]);
   generator gn465 (memory[465], 465, counter, result[465], vb[465]);
   generator gn891 (memory[891], 891, counter, result[891], vb[891]);
   generator gn768 (memory[768], 768, counter, result[768], vb[768]);
   generator gn57 (memory[57], 57, counter, result[57], vb[57]);
   generator gn718 (memory[718], 718, counter, result[718], vb[718]);
   generator gn91 (memory[91], 91, counter, result[91], vb[91]);
   generator gn764 (memory[764], 764, counter, result[764], vb[764]);
   generator gn829 (memory[829], 829, counter, result[829], vb[829]);
   generator gn892 (memory[892], 892, counter, result[892], vb[892]);
   generator gn140 (memory[140], 140, counter, result[140], vb[140]);
   generator gn133 (memory[133], 133, counter, result[133], vb[133]);
   generator gn352 (memory[352], 352, counter, result[352], vb[352]);
   generator gn262 (memory[262], 262, counter, result[262], vb[262]);
   generator gn868 (memory[868], 868, counter, result[868], vb[868]);
   generator gn296 (memory[296], 296, counter, result[296], vb[296]);
   generator gn191 (memory[191], 191, counter, result[191], vb[191]);
   generator gn652 (memory[652], 652, counter, result[652], vb[652]);
   generator gn413 (memory[413], 413, counter, result[413], vb[413]);
   generator gn437 (memory[437], 437, counter, result[437], vb[437]);
   generator gn944 (memory[944], 944, counter, result[944], vb[944]);
   generator gn694 (memory[694], 694, counter, result[694], vb[694]);
   generator gn67 (memory[67], 67, counter, result[67], vb[67]);
   generator gn509 (memory[509], 509, counter, result[509], vb[509]);
   generator gn60 (memory[60], 60, counter, result[60], vb[60]);
   generator gn806 (memory[806], 806, counter, result[806], vb[806]);
   generator gn490 (memory[490], 490, counter, result[490], vb[490]);
   generator gn155 (memory[155], 155, counter, result[155], vb[155]);
   generator gn882 (memory[882], 882, counter, result[882], vb[882]);
   generator gn427 (memory[427], 427, counter, result[427], vb[427]);
   generator gn475 (memory[475], 475, counter, result[475], vb[475]);
   generator gn319 (memory[319], 319, counter, result[319], vb[319]);
   generator gn282 (memory[282], 282, counter, result[282], vb[282]);
   generator gn820 (memory[820], 820, counter, result[820], vb[820]);
   generator gn435 (memory[435], 435, counter, result[435], vb[435]);
   generator gn314 (memory[314], 314, counter, result[314], vb[314]);
   generator gn485 (memory[485], 485, counter, result[485], vb[485]);
   generator gn252 (memory[252], 252, counter, result[252], vb[252]);
   generator gn886 (memory[886], 886, counter, result[886], vb[886]);
   generator gn880 (memory[880], 880, counter, result[880], vb[880]);
   generator gn266 (memory[266], 266, counter, result[266], vb[266]);
   generator gn644 (memory[644], 644, counter, result[644], vb[644]);
   generator gn876 (memory[876], 876, counter, result[876], vb[876]);
   generator gn206 (memory[206], 206, counter, result[206], vb[206]);
   generator gn312 (memory[312], 312, counter, result[312], vb[312]);
   generator gn628 (memory[628], 628, counter, result[628], vb[628]);
   generator gn280 (memory[280], 280, counter, result[280], vb[280]);
   generator gn970 (memory[970], 970, counter, result[970], vb[970]);
   generator gn150 (memory[150], 150, counter, result[150], vb[150]);
   generator gn630 (memory[630], 630, counter, result[630], vb[630]);
   generator gn457 (memory[457], 457, counter, result[457], vb[457]);
   generator gn163 (memory[163], 163, counter, result[163], vb[163]);
   generator gn269 (memory[269], 269, counter, result[269], vb[269]);
   generator gn24 (memory[24], 24, counter, result[24], vb[24]);
   generator gn834 (memory[834], 834, counter, result[834], vb[834]);
   generator gn862 (memory[862], 862, counter, result[862], vb[862]);
   generator gn674 (memory[674], 674, counter, result[674], vb[674]);
   generator gn87 (memory[87], 87, counter, result[87], vb[87]);
   generator gn541 (memory[541], 541, counter, result[541], vb[541]);
   generator gn146 (memory[146], 146, counter, result[146], vb[146]);
   generator gn386 (memory[386], 386, counter, result[386], vb[386]);
   generator gn419 (memory[419], 419, counter, result[419], vb[419]);
   generator gn28 (memory[28], 28, counter, result[28], vb[28]);
   generator gn612 (memory[612], 612, counter, result[612], vb[612]);
   generator gn747 (memory[747], 747, counter, result[747], vb[747]);
   generator gn129 (memory[129], 129, counter, result[129], vb[129]);
   generator gn180 (memory[180], 180, counter, result[180], vb[180]);
   generator gn741 (memory[741], 741, counter, result[741], vb[741]);
   generator gn179 (memory[179], 179, counter, result[179], vb[179]);
   generator gn523 (memory[523], 523, counter, result[523], vb[523]);
   generator gn62 (memory[62], 62, counter, result[62], vb[62]);
   generator gn430 (memory[430], 430, counter, result[430], vb[430]);
   generator gn251 (memory[251], 251, counter, result[251], vb[251]);
   generator gn479 (memory[479], 479, counter, result[479], vb[479]);
   generator gn199 (memory[199], 199, counter, result[199], vb[199]);
   generator gn478 (memory[478], 478, counter, result[478], vb[478]);
   generator gn669 (memory[669], 669, counter, result[669], vb[669]);
   generator gn460 (memory[460], 460, counter, result[460], vb[460]);
   generator gn392 (memory[392], 392, counter, result[392], vb[392]);
   generator gn662 (memory[662], 662, counter, result[662], vb[662]);
   generator gn170 (memory[170], 170, counter, result[170], vb[170]);
   generator gn425 (memory[425], 425, counter, result[425], vb[425]);
   generator gn898 (memory[898], 898, counter, result[898], vb[898]);
   generator gn870 (memory[870], 870, counter, result[870], vb[870]);
   generator gn548 (memory[548], 548, counter, result[548], vb[548]);
   generator gn581 (memory[581], 581, counter, result[581], vb[581]);
   generator gn813 (memory[813], 813, counter, result[813], vb[813]);
   generator gn388 (memory[388], 388, counter, result[388], vb[388]);
   generator gn436 (memory[436], 436, counter, result[436], vb[436]);
   generator gn245 (memory[245], 245, counter, result[245], vb[245]);
   generator gn881 (memory[881], 881, counter, result[881], vb[881]);
   generator gn167 (memory[167], 167, counter, result[167], vb[167]);
   generator gn173 (memory[173], 173, counter, result[173], vb[173]);
   generator gn442 (memory[442], 442, counter, result[442], vb[442]);
   generator gn525 (memory[525], 525, counter, result[525], vb[525]);
   generator gn363 (memory[363], 363, counter, result[363], vb[363]);
   generator gn826 (memory[826], 826, counter, result[826], vb[826]);
   generator gn211 (memory[211], 211, counter, result[211], vb[211]);
   generator gn608 (memory[608], 608, counter, result[608], vb[608]);
   generator gn914 (memory[914], 914, counter, result[914], vb[914]);
   generator gn408 (memory[408], 408, counter, result[408], vb[408]);
   generator gn186 (memory[186], 186, counter, result[186], vb[186]);
   generator gn399 (memory[399], 399, counter, result[399], vb[399]);
   generator gn507 (memory[507], 507, counter, result[507], vb[507]);
   generator gn936 (memory[936], 936, counter, result[936], vb[936]);
   generator gn422 (memory[422], 422, counter, result[422], vb[422]);
   generator gn300 (memory[300], 300, counter, result[300], vb[300]);
   generator gn302 (memory[302], 302, counter, result[302], vb[302]);
   generator gn118 (memory[118], 118, counter, result[118], vb[118]);
   generator gn209 (memory[209], 209, counter, result[209], vb[209]);
   generator gn974 (memory[974], 974, counter, result[974], vb[974]);
   generator gn879 (memory[879], 879, counter, result[879], vb[879]);
   generator gn896 (memory[896], 896, counter, result[896], vb[896]);
   generator gn993 (memory[993], 993, counter, result[993], vb[993]);
   generator gn286 (memory[286], 286, counter, result[286], vb[286]);
   generator gn654 (memory[654], 654, counter, result[654], vb[654]);
   generator gn440 (memory[440], 440, counter, result[440], vb[440]);
   generator gn107 (memory[107], 107, counter, result[107], vb[107]);
   generator gn735 (memory[735], 735, counter, result[735], vb[735]);
   generator gn250 (memory[250], 250, counter, result[250], vb[250]);
   generator gn871 (memory[871], 871, counter, result[871], vb[871]);
   generator gn976 (memory[976], 976, counter, result[976], vb[976]);
   generator gn117 (memory[117], 117, counter, result[117], vb[117]);
   generator gn356 (memory[356], 356, counter, result[356], vb[356]);
   generator gn92 (memory[92], 92, counter, result[92], vb[92]);
   generator gn505 (memory[505], 505, counter, result[505], vb[505]);
   generator gn783 (memory[783], 783, counter, result[783], vb[783]);
   generator gn809 (memory[809], 809, counter, result[809], vb[809]);
   generator gn246 (memory[246], 246, counter, result[246], vb[246]);
   generator gn382 (memory[382], 382, counter, result[382], vb[382]);
   generator gn589 (memory[589], 589, counter, result[589], vb[589]);
   generator gn994 (memory[994], 994, counter, result[994], vb[994]);
   generator gn304 (memory[304], 304, counter, result[304], vb[304]);
   generator gn760 (memory[760], 760, counter, result[760], vb[760]);
   generator gn78 (memory[78], 78, counter, result[78], vb[78]);
   generator gn410 (memory[410], 410, counter, result[410], vb[410]);
   generator gn390 (memory[390], 390, counter, result[390], vb[390]);
   generator gn48 (memory[48], 48, counter, result[48], vb[48]);
   generator gn89 (memory[89], 89, counter, result[89], vb[89]);
   generator gn201 (memory[201], 201, counter, result[201], vb[201]);
   generator gn869 (memory[869], 869, counter, result[869], vb[869]);
   generator gn831 (memory[831], 831, counter, result[831], vb[831]);
   generator gn894 (memory[894], 894, counter, result[894], vb[894]);
   generator gn149 (memory[149], 149, counter, result[149], vb[149]);
   generator gn971 (memory[971], 971, counter, result[971], vb[971]);
   generator gn865 (memory[865], 865, counter, result[865], vb[865]);
   generator gn928 (memory[928], 928, counter, result[928], vb[928]);
   generator gn369 (memory[369], 369, counter, result[369], vb[369]);
   generator gn52 (memory[52], 52, counter, result[52], vb[52]);
   generator gn6 (memory[6], 6, counter, result[6], vb[6]);
   generator gn565 (memory[565], 565, counter, result[565], vb[565]);
   generator gn979 (memory[979], 979, counter, result[979], vb[979]);
   generator gn743 (memory[743], 743, counter, result[743], vb[743]);
   generator gn177 (memory[177], 177, counter, result[177], vb[177]);
   generator gn655 (memory[655], 655, counter, result[655], vb[655]);
   generator gn812 (memory[812], 812, counter, result[812], vb[812]);
   generator gn277 (memory[277], 277, counter, result[277], vb[277]);
   generator gn846 (memory[846], 846, counter, result[846], vb[846]);
   generator gn341 (memory[341], 341, counter, result[341], vb[341]);
   generator gn853 (memory[853], 853, counter, result[853], vb[853]);
   generator gn819 (memory[819], 819, counter, result[819], vb[819]);
   generator gn945 (memory[945], 945, counter, result[945], vb[945]);
   generator gn1017 (memory[1017], 1017, counter, result[1017], vb[1017]);
   generator gn591 (memory[591], 591, counter, result[591], vb[591]);
   generator gn194 (memory[194], 194, counter, result[194], vb[194]);
   generator gn653 (memory[653], 653, counter, result[653], vb[653]);
   generator gn114 (memory[114], 114, counter, result[114], vb[114]);
   generator gn313 (memory[313], 313, counter, result[313], vb[313]);
   generator gn506 (memory[506], 506, counter, result[506], vb[506]);
   generator gn21 (memory[21], 21, counter, result[21], vb[21]);
   generator gn351 (memory[351], 351, counter, result[351], vb[351]);
   generator gn486 (memory[486], 486, counter, result[486], vb[486]);
   generator gn330 (memory[330], 330, counter, result[330], vb[330]);
   generator gn875 (memory[875], 875, counter, result[875], vb[875]);
   generator gn139 (memory[139], 139, counter, result[139], vb[139]);
   generator gn1011 (memory[1011], 1011, counter, result[1011], vb[1011]);
   generator gn877 (memory[877], 877, counter, result[877], vb[877]);
   generator gn458 (memory[458], 458, counter, result[458], vb[458]);
   generator gn751 (memory[751], 751, counter, result[751], vb[751]);
   generator gn217 (memory[217], 217, counter, result[217], vb[217]);
   generator gn42 (memory[42], 42, counter, result[42], vb[42]);
   generator gn930 (memory[930], 930, counter, result[930], vb[930]);
   generator gn641 (memory[641], 641, counter, result[641], vb[641]);
   generator gn58 (memory[58], 58, counter, result[58], vb[58]);
   generator gn342 (memory[342], 342, counter, result[342], vb[342]);
   generator gn165 (memory[165], 165, counter, result[165], vb[165]);
   generator gn750 (memory[750], 750, counter, result[750], vb[750]);
   generator gn258 (memory[258], 258, counter, result[258], vb[258]);
   generator gn948 (memory[948], 948, counter, result[948], vb[948]);
   generator gn961 (memory[961], 961, counter, result[961], vb[961]);
   generator gn682 (memory[682], 682, counter, result[682], vb[682]);
   generator gn1007 (memory[1007], 1007, counter, result[1007], vb[1007]);
   generator gn265 (memory[265], 265, counter, result[265], vb[265]);
   generator gn709 (memory[709], 709, counter, result[709], vb[709]);
   generator gn978 (memory[978], 978, counter, result[978], vb[978]);
   generator gn726 (memory[726], 726, counter, result[726], vb[726]);
   generator gn497 (memory[497], 497, counter, result[497], vb[497]);
   generator gn695 (memory[695], 695, counter, result[695], vb[695]);
   generator gn355 (memory[355], 355, counter, result[355], vb[355]);
   generator gn510 (memory[510], 510, counter, result[510], vb[510]);
   generator gn511 (memory[511], 511, counter, result[511], vb[511]);
   generator gn987 (memory[987], 987, counter, result[987], vb[987]);
   generator gn555 (memory[555], 555, counter, result[555], vb[555]);
   generator gn714 (memory[714], 714, counter, result[714], vb[714]);
   generator gn10 (memory[10], 10, counter, result[10], vb[10]);
   generator gn666 (memory[666], 666, counter, result[666], vb[666]);
   generator gn72 (memory[72], 72, counter, result[72], vb[72]);
   generator gn320 (memory[320], 320, counter, result[320], vb[320]);
   generator gn278 (memory[278], 278, counter, result[278], vb[278]);
   generator gn379 (memory[379], 379, counter, result[379], vb[379]);
   generator gn549 (memory[549], 549, counter, result[549], vb[549]);
   generator gn339 (memory[339], 339, counter, result[339], vb[339]);
   generator gn7 (memory[7], 7, counter, result[7], vb[7]);
   generator gn53 (memory[53], 53, counter, result[53], vb[53]);
   generator gn164 (memory[164], 164, counter, result[164], vb[164]);
   generator gn321 (memory[321], 321, counter, result[321], vb[321]);
   generator gn401 (memory[401], 401, counter, result[401], vb[401]);
   generator gn242 (memory[242], 242, counter, result[242], vb[242]);
   generator gn71 (memory[71], 71, counter, result[71], vb[71]);
   generator gn285 (memory[285], 285, counter, result[285], vb[285]);
   generator gn272 (memory[272], 272, counter, result[272], vb[272]);
   generator gn965 (memory[965], 965, counter, result[965], vb[965]);
   generator gn367 (memory[367], 367, counter, result[367], vb[367]);
   generator gn958 (memory[958], 958, counter, result[958], vb[958]);
   generator gn611 (memory[611], 611, counter, result[611], vb[611]);
   generator gn1016 (memory[1016], 1016, counter, result[1016], vb[1016]);
   generator gn704 (memory[704], 704, counter, result[704], vb[704]);
   generator gn215 (memory[215], 215, counter, result[215], vb[215]);
   generator gn539 (memory[539], 539, counter, result[539], vb[539]);
   generator gn32 (memory[32], 32, counter, result[32], vb[32]);
   generator gn765 (memory[765], 765, counter, result[765], vb[765]);
   generator gn706 (memory[706], 706, counter, result[706], vb[706]);
   generator gn545 (memory[545], 545, counter, result[545], vb[545]);
   generator gn723 (memory[723], 723, counter, result[723], vb[723]);
   generator gn403 (memory[403], 403, counter, result[403], vb[403]);
   generator gn103 (memory[103], 103, counter, result[103], vb[103]);
   generator gn687 (memory[687], 687, counter, result[687], vb[687]);
   generator gn185 (memory[185], 185, counter, result[185], vb[185]);
   generator gn609 (memory[609], 609, counter, result[609], vb[609]);
   generator gn696 (memory[696], 696, counter, result[696], vb[696]);
   generator gn623 (memory[623], 623, counter, result[623], vb[623]);
   generator gn152 (memory[152], 152, counter, result[152], vb[152]);
   generator gn239 (memory[239], 239, counter, result[239], vb[239]);
   generator gn901 (memory[901], 901, counter, result[901], vb[901]);
   generator gn452 (memory[452], 452, counter, result[452], vb[452]);
   generator gn632 (memory[632], 632, counter, result[632], vb[632]);
   generator gn256 (memory[256], 256, counter, result[256], vb[256]);
   generator gn4 (memory[4], 4, counter, result[4], vb[4]);
   generator gn665 (memory[665], 665, counter, result[665], vb[665]);
   generator gn79 (memory[79], 79, counter, result[79], vb[79]);
   generator gn782 (memory[782], 782, counter, result[782], vb[782]);
   generator gn8 (memory[8], 8, counter, result[8], vb[8]);
   generator gn415 (memory[415], 415, counter, result[415], vb[415]);
   generator gn450 (memory[450], 450, counter, result[450], vb[450]);
   generator gn270 (memory[270], 270, counter, result[270], vb[270]);
   generator gn168 (memory[168], 168, counter, result[168], vb[168]);
   generator gn855 (memory[855], 855, counter, result[855], vb[855]);
   generator gn660 (memory[660], 660, counter, result[660], vb[660]);
   generator gn358 (memory[358], 358, counter, result[358], vb[358]);
   generator gn333 (memory[333], 333, counter, result[333], vb[333]);
   generator gn999 (memory[999], 999, counter, result[999], vb[999]);
   generator gn421 (memory[421], 421, counter, result[421], vb[421]);
   generator gn253 (memory[253], 253, counter, result[253], vb[253]);
   generator gn959 (memory[959], 959, counter, result[959], vb[959]);
   generator gn963 (memory[963], 963, counter, result[963], vb[963]);
   generator gn106 (memory[106], 106, counter, result[106], vb[106]);
   generator gn997 (memory[997], 997, counter, result[997], vb[997]);
   generator gn407 (memory[407], 407, counter, result[407], vb[407]);
   generator gn583 (memory[583], 583, counter, result[583], vb[583]);
   generator gn85 (memory[85], 85, counter, result[85], vb[85]);
   generator gn553 (memory[553], 553, counter, result[553], vb[553]);
   generator gn836 (memory[836], 836, counter, result[836], vb[836]);
   generator gn827 (memory[827], 827, counter, result[827], vb[827]);
   generator gn396 (memory[396], 396, counter, result[396], vb[396]);
   generator gn197 (memory[197], 197, counter, result[197], vb[197]);
   generator gn626 (memory[626], 626, counter, result[626], vb[626]);
   generator gn573 (memory[573], 573, counter, result[573], vb[573]);
   generator gn190 (memory[190], 190, counter, result[190], vb[190]);
   generator gn88 (memory[88], 88, counter, result[88], vb[88]);
   generator gn736 (memory[736], 736, counter, result[736], vb[736]);
   generator gn417 (memory[417], 417, counter, result[417], vb[417]);
   generator gn134 (memory[134], 134, counter, result[134], vb[134]);
   generator gn283 (memory[283], 283, counter, result[283], vb[283]);
   generator gn132 (memory[132], 132, counter, result[132], vb[132]);
   generator gn814 (memory[814], 814, counter, result[814], vb[814]);
   generator gn552 (memory[552], 552, counter, result[552], vb[552]);
   generator gn82 (memory[82], 82, counter, result[82], vb[82]);
   generator gn818 (memory[818], 818, counter, result[818], vb[818]);
   generator gn236 (memory[236], 236, counter, result[236], vb[236]);
   generator gn196 (memory[196], 196, counter, result[196], vb[196]);
   generator gn224 (memory[224], 224, counter, result[224], vb[224]);
   generator gn796 (memory[796], 796, counter, result[796], vb[796]);
   generator gn1015 (memory[1015], 1015, counter, result[1015], vb[1015]);
   generator gn5 (memory[5], 5, counter, result[5], vb[5]);
   generator gn592 (memory[592], 592, counter, result[592], vb[592]);
   generator gn689 (memory[689], 689, counter, result[689], vb[689]);
   generator gn1006 (memory[1006], 1006, counter, result[1006], vb[1006]);
   generator gn471 (memory[471], 471, counter, result[471], vb[471]);
   generator gn366 (memory[366], 366, counter, result[366], vb[366]);
   generator gn301 (memory[301], 301, counter, result[301], vb[301]);
   generator gn739 (memory[739], 739, counter, result[739], vb[739]);
   generator gn745 (memory[745], 745, counter, result[745], vb[745]);
   generator gn848 (memory[848], 848, counter, result[848], vb[848]);
   generator gn193 (memory[193], 193, counter, result[193], vb[193]);
   generator gn952 (memory[952], 952, counter, result[952], vb[952]);
   generator gn461 (memory[461], 461, counter, result[461], vb[461]);
   generator gn807 (memory[807], 807, counter, result[807], vb[807]);
   generator gn254 (memory[254], 254, counter, result[254], vb[254]);
   generator gn544 (memory[544], 544, counter, result[544], vb[544]);
   generator gn964 (memory[964], 964, counter, result[964], vb[964]);
   generator gn614 (memory[614], 614, counter, result[614], vb[614]);
   generator gn77 (memory[77], 77, counter, result[77], vb[77]);
   generator gn443 (memory[443], 443, counter, result[443], vb[443]);
   generator gn561 (memory[561], 561, counter, result[561], vb[561]);
   generator gn64 (memory[64], 64, counter, result[64], vb[64]);
   generator gn940 (memory[940], 940, counter, result[940], vb[940]);
   generator gn214 (memory[214], 214, counter, result[214], vb[214]);
   generator gn378 (memory[378], 378, counter, result[378], vb[378]);
   generator gn788 (memory[788], 788, counter, result[788], vb[788]);
   generator gn610 (memory[610], 610, counter, result[610], vb[610]);
   generator gn348 (memory[348], 348, counter, result[348], vb[348]);
   generator gn1003 (memory[1003], 1003, counter, result[1003], vb[1003]);
   generator gn697 (memory[697], 697, counter, result[697], vb[697]);
   generator gn426 (memory[426], 426, counter, result[426], vb[426]);
   generator gn946 (memory[946], 946, counter, result[946], vb[946]);
   generator gn18 (memory[18], 18, counter, result[18], vb[18]);
   generator gn350 (memory[350], 350, counter, result[350], vb[350]);
   generator gn607 (memory[607], 607, counter, result[607], vb[607]);
   generator gn445 (memory[445], 445, counter, result[445], vb[445]);
   generator gn540 (memory[540], 540, counter, result[540], vb[540]);
   generator gn373 (memory[373], 373, counter, result[373], vb[373]);
   generator gn969 (memory[969], 969, counter, result[969], vb[969]);
   generator gn922 (memory[922], 922, counter, result[922], vb[922]);
   generator gn1022 (memory[1022], 1022, counter, result[1022], vb[1022]);
   generator gn377 (memory[377], 377, counter, result[377], vb[377]);
   generator gn240 (memory[240], 240, counter, result[240], vb[240]);
   generator gn778 (memory[778], 778, counter, result[778], vb[778]);
   generator gn859 (memory[859], 859, counter, result[859], vb[859]);
   generator gn520 (memory[520], 520, counter, result[520], vb[520]);
   generator gn574 (memory[574], 574, counter, result[574], vb[574]);
   generator gn636 (memory[636], 636, counter, result[636], vb[636]);
   generator gn44 (memory[44], 44, counter, result[44], vb[44]);
   generator gn531 (memory[531], 531, counter, result[531], vb[531]);
   generator gn332 (memory[332], 332, counter, result[332], vb[332]);
   generator gn261 (memory[261], 261, counter, result[261], vb[261]);
   generator gn960 (memory[960], 960, counter, result[960], vb[960]);
   generator gn564 (memory[564], 564, counter, result[564], vb[564]);
   generator gn911 (memory[911], 911, counter, result[911], vb[911]);
   generator gn447 (memory[447], 447, counter, result[447], vb[447]);
   generator gn762 (memory[762], 762, counter, result[762], vb[762]);
   generator gn594 (memory[594], 594, counter, result[594], vb[594]);
   generator gn558 (memory[558], 558, counter, result[558], vb[558]);
   generator gn257 (memory[257], 257, counter, result[257], vb[257]);
   generator gn448 (memory[448], 448, counter, result[448], vb[448]);
   generator gn716 (memory[716], 716, counter, result[716], vb[716]);
   generator gn234 (memory[234], 234, counter, result[234], vb[234]);
   generator gn222 (memory[222], 222, counter, result[222], vb[222]);
   generator gn477 (memory[477], 477, counter, result[477], vb[477]);
   generator gn754 (memory[754], 754, counter, result[754], vb[754]);
   generator gn147 (memory[147], 147, counter, result[147], vb[147]);
   generator gn213 (memory[213], 213, counter, result[213], vb[213]);
   generator gn973 (memory[973], 973, counter, result[973], vb[973]);
   generator gn667 (memory[667], 667, counter, result[667], vb[667]);
   generator gn512 (memory[512], 512, counter, result[512], vb[512]);
   generator gn264 (memory[264], 264, counter, result[264], vb[264]);
   generator gn530 (memory[530], 530, counter, result[530], vb[530]);
   generator gn65 (memory[65], 65, counter, result[65], vb[65]);
   generator gn658 (memory[658], 658, counter, result[658], vb[658]);
   generator gn128 (memory[128], 128, counter, result[128], vb[128]);
   generator gn986 (memory[986], 986, counter, result[986], vb[986]);
   generator gn126 (memory[126], 126, counter, result[126], vb[126]);
   generator gn670 (memory[670], 670, counter, result[670], vb[670]);
   generator gn800 (memory[800], 800, counter, result[800], vb[800]);
   generator gn238 (memory[238], 238, counter, result[238], vb[238]);
   generator gn353 (memory[353], 353, counter, result[353], vb[353]);
   generator gn563 (memory[563], 563, counter, result[563], vb[563]);
   generator gn294 (memory[294], 294, counter, result[294], vb[294]);
   generator gn954 (memory[954], 954, counter, result[954], vb[954]);
   generator gn428 (memory[428], 428, counter, result[428], vb[428]);
   generator gn488 (memory[488], 488, counter, result[488], vb[488]);
   generator gn235 (memory[235], 235, counter, result[235], vb[235]);
   generator gn989 (memory[989], 989, counter, result[989], vb[989]);
   generator gn801 (memory[801], 801, counter, result[801], vb[801]);
   generator gn281 (memory[281], 281, counter, result[281], vb[281]);
   generator gn514 (memory[514], 514, counter, result[514], vb[514]);
   generator gn375 (memory[375], 375, counter, result[375], vb[375]);
   generator gn631 (memory[631], 631, counter, result[631], vb[631]);
   generator gn534 (memory[534], 534, counter, result[534], vb[534]);
   generator gn210 (memory[210], 210, counter, result[210], vb[210]);
   generator gn385 (memory[385], 385, counter, result[385], vb[385]);
   generator gn772 (memory[772], 772, counter, result[772], vb[772]);
   generator gn141 (memory[141], 141, counter, result[141], vb[141]);
   generator gn459 (memory[459], 459, counter, result[459], vb[459]);
   generator gn982 (memory[982], 982, counter, result[982], vb[982]);
   generator gn947 (memory[947], 947, counter, result[947], vb[947]);
   generator gn484 (memory[484], 484, counter, result[484], vb[484]);
   generator gn61 (memory[61], 61, counter, result[61], vb[61]);
   generator gn748 (memory[748], 748, counter, result[748], vb[748]);
   generator gn516 (memory[516], 516, counter, result[516], vb[516]);
   generator gn912 (memory[912], 912, counter, result[912], vb[912]);
   generator gn41 (memory[41], 41, counter, result[41], vb[41]);
   generator gn416 (memory[416], 416, counter, result[416], vb[416]);
   generator gn677 (memory[677], 677, counter, result[677], vb[677]);
   generator gn36 (memory[36], 36, counter, result[36], vb[36]);
   generator gn221 (memory[221], 221, counter, result[221], vb[221]);
   generator gn538 (memory[538], 538, counter, result[538], vb[538]);
   generator gn481 (memory[481], 481, counter, result[481], vb[481]);
   generator gn145 (memory[145], 145, counter, result[145], vb[145]);
   generator gn500 (memory[500], 500, counter, result[500], vb[500]);
   generator gn212 (memory[212], 212, counter, result[212], vb[212]);
   generator gn502 (memory[502], 502, counter, result[502], vb[502]);
   generator gn863 (memory[863], 863, counter, result[863], vb[863]);
   generator gn618 (memory[618], 618, counter, result[618], vb[618]);
   generator gn576 (memory[576], 576, counter, result[576], vb[576]);
   generator gn551 (memory[551], 551, counter, result[551], vb[551]);
   generator gn556 (memory[556], 556, counter, result[556], vb[556]);
   generator gn409 (memory[409], 409, counter, result[409], vb[409]);
   generator gn306 (memory[306], 306, counter, result[306], vb[306]);
   generator gn532 (memory[532], 532, counter, result[532], vb[532]);
   generator gn830 (memory[830], 830, counter, result[830], vb[830]);
   generator gn799 (memory[799], 799, counter, result[799], vb[799]);
   generator gn51 (memory[51], 51, counter, result[51], vb[51]);
   generator gn861 (memory[861], 861, counter, result[861], vb[861]);
   generator gn643 (memory[643], 643, counter, result[643], vb[643]);
   generator gn749 (memory[749], 749, counter, result[749], vb[749]);
   generator gn287 (memory[287], 287, counter, result[287], vb[287]);
   generator gn371 (memory[371], 371, counter, result[371], vb[371]);
   generator gn821 (memory[821], 821, counter, result[821], vb[821]);
   generator gn795 (memory[795], 795, counter, result[795], vb[795]);
   generator gn937 (memory[937], 937, counter, result[937], vb[937]);
   generator gn455 (memory[455], 455, counter, result[455], vb[455]);
   generator gn404 (memory[404], 404, counter, result[404], vb[404]);
   generator gn776 (memory[776], 776, counter, result[776], vb[776]);
   generator gn169 (memory[169], 169, counter, result[169], vb[169]);
   generator gn166 (memory[166], 166, counter, result[166], vb[166]);
   generator gn663 (memory[663], 663, counter, result[663], vb[663]);
   generator gn151 (memory[151], 151, counter, result[151], vb[151]);
   generator gn810 (memory[810], 810, counter, result[810], vb[810]);
   generator gn112 (memory[112], 112, counter, result[112], vb[112]);
   generator gn244 (memory[244], 244, counter, result[244], vb[244]);
   generator gn39 (memory[39], 39, counter, result[39], vb[39]);
   generator gn192 (memory[192], 192, counter, result[192], vb[192]);
   generator gn70 (memory[70], 70, counter, result[70], vb[70]);
   generator gn393 (memory[393], 393, counter, result[393], vb[393]);
   generator gn580 (memory[580], 580, counter, result[580], vb[580]);
   generator gn887 (memory[887], 887, counter, result[887], vb[887]);
   generator gn910 (memory[910], 910, counter, result[910], vb[910]);
   generator gn890 (memory[890], 890, counter, result[890], vb[890]);
   generator gn131 (memory[131], 131, counter, result[131], vb[131]);
   generator gn324 (memory[324], 324, counter, result[324], vb[324]);
   generator gn136 (memory[136], 136, counter, result[136], vb[136]);
   generator gn411 (memory[411], 411, counter, result[411], vb[411]);
   generator gn688 (memory[688], 688, counter, result[688], vb[688]);
   generator gn983 (memory[983], 983, counter, result[983], vb[983]);
   generator gn307 (memory[307], 307, counter, result[307], vb[307]);
   generator gn524 (memory[524], 524, counter, result[524], vb[524]);
   generator gn19 (memory[19], 19, counter, result[19], vb[19]);
   generator gn543 (memory[543], 543, counter, result[543], vb[543]);
   generator gn1009 (memory[1009], 1009, counter, result[1009], vb[1009]);
   generator gn815 (memory[815], 815, counter, result[815], vb[815]);
   generator gn233 (memory[233], 233, counter, result[233], vb[233]);
   generator gn496 (memory[496], 496, counter, result[496], vb[496]);
   generator gn906 (memory[906], 906, counter, result[906], vb[906]);
   generator gn752 (memory[752], 752, counter, result[752], vb[752]);
   generator gn816 (memory[816], 816, counter, result[816], vb[816]);
   generator gn738 (memory[738], 738, counter, result[738], vb[738]);
   generator gn95 (memory[95], 95, counter, result[95], vb[95]);
   generator gn582 (memory[582], 582, counter, result[582], vb[582]);
   generator gn494 (memory[494], 494, counter, result[494], vb[494]);
   generator gn640 (memory[640], 640, counter, result[640], vb[640]);
   generator gn872 (memory[872], 872, counter, result[872], vb[872]);
   generator gn924 (memory[924], 924, counter, result[924], vb[924]);
   generator gn761 (memory[761], 761, counter, result[761], vb[761]);
   generator gn55 (memory[55], 55, counter, result[55], vb[55]);
   generator gn116 (memory[116], 116, counter, result[116], vb[116]);
   generator gn47 (memory[47], 47, counter, result[47], vb[47]);
   generator gn518 (memory[518], 518, counter, result[518], vb[518]);
   generator gn259 (memory[259], 259, counter, result[259], vb[259]);
   generator gn664 (memory[664], 664, counter, result[664], vb[664]);
   generator gn980 (memory[980], 980, counter, result[980], vb[980]);
   generator gn115 (memory[115], 115, counter, result[115], vb[115]);
   generator gn586 (memory[586], 586, counter, result[586], vb[586]);
   generator gn988 (memory[988], 988, counter, result[988], vb[988]);
   generator gn587 (memory[587], 587, counter, result[587], vb[587]);
   generator gn878 (memory[878], 878, counter, result[878], vb[878]);
   generator gn647 (memory[647], 647, counter, result[647], vb[647]);
   generator gn205 (memory[205], 205, counter, result[205], vb[205]);
   generator gn480 (memory[480], 480, counter, result[480], vb[480]);
   generator gn925 (memory[925], 925, counter, result[925], vb[925]);
   generator gn20 (memory[20], 20, counter, result[20], vb[20]);
   generator gn672 (memory[672], 672, counter, result[672], vb[672]);
   generator gn727 (memory[727], 727, counter, result[727], vb[727]);
   generator gn559 (memory[559], 559, counter, result[559], vb[559]);
   generator gn123 (memory[123], 123, counter, result[123], vb[123]);
   generator gn446 (memory[446], 446, counter, result[446], vb[446]);
   generator gn176 (memory[176], 176, counter, result[176], vb[176]);
   generator gn710 (memory[710], 710, counter, result[710], vb[710]);
   generator gn83 (memory[83], 83, counter, result[83], vb[83]);
   generator gn918 (memory[918], 918, counter, result[918], vb[918]);
   generator gn429 (memory[429], 429, counter, result[429], vb[429]);
   generator gn803 (memory[803], 803, counter, result[803], vb[803]);
   generator gn966 (memory[966], 966, counter, result[966], vb[966]);
   generator gn308 (memory[308], 308, counter, result[308], vb[308]);
   
   initial begin
       counter = 0;
       memory[323] = 144'hfe354ea23e90ba0dd0024f530da99bf732fc;
       memory[257] = 144'h16ca4d36dea8fa09dfd003dcb53a3a43888f;
       memory[427] = 144'ha93602f4716f1a0b7bf316643736710003a5;
       memory[336] = 144'h728c67a98e5efa224ab23306a406ca2a0cbd;
       memory[143] = 144'hea300a26b3d9602754f95d6539f0af8ba02b;
       memory[273] = 144'h71af463e7ee1632716fab30266c4db76a118;
       memory[389] = 144'hd9ec4f723c22ab4cd32d8e6320567244f420;
       memory[523] = 144'hf87d064a9213c26f55e6e9b6d28491b94726;
       memory[147] = 144'ha29f04a75007652bd2d8903bcf684c4e1ec7;
       memory[179] = 144'h932303f2d071010fcc40ebe7a2d3e37d9772;
       memory[146] = 144'heba62f063070fc00522ac15a634d68b5d431;
       memory[516] = 144'h470262162ea498085319964a9746ab5f47d2;
       memory[385] = 144'ha68d45451ebdea20f8385073ded52abee211;
       memory[375] = 144'hb5414d04fe4abc2fa3684a34afed96e0405b;
       memory[376] = 144'h46436bc9ce236304ed4869c30c46947ec1b4;
       memory[43] = 144'ha5d104437058b72cc7bac57c1e816ef76e9e;
       memory[378] = 144'h8e866fc35ed41b085018f9089902c3393d32;
       memory[34] = 144'hde5f24a430349227016078e0812852604ff7;
       memory[99] = 144'haeff09f8525ff1441e7f10a3a2e86156580d;
       memory[580] = 144'h268766975f797e2d95213ae4a1cc7cdd6bd9;
       memory[114] = 144'h78152c15d270b76f909ff7e9b50cdda5bcae;
       memory[117] = 144'hf17040171fae5668ee46dce21c92e77120a8;
       memory[424] = 144'hacd22e8c01de9e269e903d50818da52ce1fc;
       memory[563] = 144'hcff74d5b5fa5ae052561839e84d265a347a8;
       memory[540] = 144'h48496117ade721083e8809612a6882f49dfa;
       memory[123] = 144'hf0b0432e5ea82e63d95474e710a195bad2e5;
       memory[120] = 144'hb7da611d6d6acc4e0e44a8ac28f9eaba5a20;
       memory[402] = 144'haa11622cdc582428f930b3c9c573525a60bb;
       memory[617] = 144'h3d4b47923d770625f189e8360c8eaa857a26;
       memory[425] = 144'hb51102bc6131930423402df3ad3827d2c4c5;
       memory[28] = 144'h1ab9290b70515a249ee0976b10e99e30c4a3;
       memory[254] = 144'h8ac629c4b325ed2e8b23dcb0e6c5af0b7d29;
       memory[537] = 144'h770a0b63424a2d6487e6a7068e5357d41403;
       memory[49] = 144'h246c4873ef47fb654595a4f5d7779b5d075c;
       memory[352] = 144'h53f267ff3e17dc0a12c89555c74f69bfff07;
       memory[217] = 144'hb7d207b243cc026766566b1ba8eb6bda3dca;
       memory[335] = 144'h15ad4e35de82520d7ec28c558de44f74f472;
       memory[448] = 144'h9da92025d265c9405a46970c764de6289d40;
       memory[32] = 144'h501d2868a0ae3c27f6808e39de49056483cd;
       memory[108] = 144'hd1026e9b0f2a21299d726330ea7ecac74100;
       memory[530] = 144'h802d6307efcf9a4fd1f56c7f49e62835569e;
       memory[349] = 144'he0744c503e2cb60ca142a6087115957190da;
       memory[247] = 144'h840c0533c0786c04226377be352314288d4b;
       memory[446] = 144'hc056223101c492431b941879527b0bd3fedf;
       memory[276] = 144'h0cc963c98eb9ed0f40ca8938ef41e58b980c;
       memory[215] = 144'hb0fc0e64d079d829a079f9562f3dd6545edc;
       memory[193] = 144'hc41a4edbbe12ad04dcd36d416570273a4ccb;
       memory[483] = 144'h45cb4cc88db44702c751a84ab98f42f3307e;
       memory[66] = 144'h80f92a2c2273c0007fa8d8be7b1784c77f25;
       memory[209] = 144'haf1f4b63fcd96923b78a62086d7871820100;
       memory[304] = 144'h63346e9b1e64df06d458fe612978317e1706;
       memory[347] = 144'hc5c149e84e14ed06eea2a74faad57cfd3bf1;
       memory[188] = 144'h1b676dfa8c1e7764d3ed7f3fe309fa379581;
       memory[110] = 144'h8a9e63cabf551226e7823a52c132777ddecb;
       memory[167] = 144'h18b4091033b79a0ee02390fa280b12a2ddb4;
       memory[576] = 144'ha7596ab73f6eb5296f0196eea016b4864533;
       memory[536] = 144'hdc5820cf029387407435ec5970ff05798c19;
       memory[194] = 144'h15dc6c1cae68570c6ee9f620d99361056cce;
       memory[340] = 144'h8dbc6cdf2e8c132fffd292f5a983a5348e91;
       memory[400] = 144'h24d9291be1dbc52ebaf03b9833b1d91f0999;
       memory[239] = 144'h25830f81c217ab0da7819d42af58e00aac38;
       memory[52] = 144'hcdf92aa0e090b84d8c77f82c3e0c657f101f;
       memory[241] = 144'hc3de040e6236ed0ebdc1ea583a81e51b2417;
       memory[359] = 144'h91914e4c2e47fa24e7f8d78dab1cc30f202a;
       memory[139] = 144'ha7900f2273e94922e29a1af375d2cefd64b3;
       memory[418] = 144'h2dfe61668c4f1326d3100dbbffe2734d3813;
       memory[317] = 144'hb76449a0fe4ec00e0a42da2aec9c65638aa8;
       memory[259] = 144'hbe974d173eca9104ce20c9d9d5f5c6eeab59;
       memory[492] = 144'h5ed220e9b34cca61f94d8229f196d783b0ed;
       memory[468] = 144'h66eb685b9c4f8e220103ec47f1f80d970432;
       memory[272] = 144'hdfc36e5dcebd4102d6cad9479deabf6eb721;
       memory[311] = 144'hc577418c7e7c760a580285619294ee6441aa;
       memory[7] = 144'hfba2033680b29d033a9018c0608e8cbdcf01;
       memory[565] = 144'h365046741f38dd074e01b8576a9c0ee80a97;
       memory[70] = 144'h6e082c01b22bf40f41a86942dded67074245;
       memory[353] = 144'h084e444f4eef5d245d184ca8ce65ab0d64bf;
       memory[77] = 144'h1015093992719e0cfd021581a6b9ad3c0634;
       memory[102] = 144'hb8c62d0822648669f55f4fd812c8e63b518e;
       memory[256] = 144'hecd568238ef2d629cda34113b11c5be1988d;
       memory[303] = 144'hed5a40b66e9ac72a13f8374c243de40b39de;
       memory[369] = 144'h3b324e3d0eed76296c28599394c2d74740e7;
       memory[297] = 144'h768249b00e3d4e22ae28171bc62e35979ec0;
       memory[187] = 144'h2e774fee2cf7254dbd3fcd55ca170525d1b4;
       memory[228] = 144'he4326a926dd81a4bdc87ff197ffd19594eea;
       memory[514] = 144'h87de6db7de578603e1e9b7b09eaadfad9be5;
       memory[326] = 144'hd834610cdeafbd20efd2c955550484d4868b;
       memory[542] = 144'h00b264a50fbd950c91c8f51b3c011a2aa1cf;
       memory[208] = 144'h62dd6db9cc7cf607c0ba2a91501d24089f92;
       memory[95] = 144'hb15b0399e257464bf64fd15ec7010e2110f9;
       memory[249] = 144'h7da507bca02c4e0a1a83408647870078f06d;
       memory[332] = 144'hf5eb66a54ea3be2b0062ed02acef9e6c86ef;
       memory[510] = 144'hba892f6583317d416017de9a64e46e826af1;
       memory[196] = 144'h40ad647cad6a5e4319362df89b482e3cd94a;
       memory[505] = 144'h29680a4b20c607436e4d7306408a708d5afe;
       memory[162] = 144'h6d492a3ee322ee20ec60b2dce3bcb06d6eae;
       memory[320] = 144'hb2d361b32e06d8230b72a5082729e9d91efa;
       memory[112] = 144'hb3e66150efd8d72e23d2df9fb67fc83e10ba;
       memory[287] = 144'hc79347e3be2a4c204abad1ea7fe6a5f2c562;
       memory[136] = 144'h46e92de43282080a6599c1c032762516ad7c;
       memory[89] = 144'h11f307a6b1b56d4f94dc7290b4fe71b78493;
       memory[230] = 144'h374e6329cd36d44ba3e5c96517b5df99d3c5;
       memory[291] = 144'h06ea41fb5c4dfe25d2aa480dbcb2e27cc111;
       memory[172] = 144'h936c23c5d03b3e2040900127899c95fc6b1c;
       memory[473] = 144'h106d46990eb9c50944b3f52e5473fb84e5bc;
       memory[313] = 144'he3724b278ebc4e0da8021d40e0fee9c3dfea;
       memory[526] = 144'hf3936ffc8dfe910315b8615aacd16cfffdfb;
       memory[229] = 144'h921a4a09fda3036ad687189271d12c4786aa;
       memory[177] = 144'hd565015c803ae1093ee34b7b7189be130aab;
       memory[319] = 144'he34c42628e7639068af248cafa9f61e608e5;
       memory[363] = 144'h6d1147871ecca720a148479032bfb470c150;
       memory[549] = 144'h8363468c9fdbd40659c1bfc0039b7d86ac18;
       memory[608] = 144'h14c36b8b4d227d01a8799826f27cdcd3ff74;
       memory[600] = 144'h1d576fed2d234c095ef95ff9b0d90392b2d0;
       memory[581] = 144'h432b48eddf68020620e3a85623865878099a;
       memory[88] = 144'h098c2ef3014d506bc5fcc3b54eb3fd6a4421;
       memory[96] = 144'hd30a6480cf1e1224e0e2b3339e9e4137ed03;
       memory[295] = 144'h83f64fb30c4da22373a84d667082f48c35c0;
       memory[131] = 144'haaad0ee6c18d372eba2a964cdb22927045ff;
       memory[307] = 144'h7a26486c1ecd842ee8d80d92bd3a6e1f3cb7;
       memory[460] = 144'h32c725c1516d4c4988e48d9f24b0c7706ece;
       memory[439] = 144'h4cc40a5e50cca32450f980d5688100f10162;
       memory[588] = 144'hbd3d60b1cda8ca0a77392c3ac920386eca64;
       memory[545] = 144'h695e412cefee870494019ad41befe4138a2b;
       memory[480] = 144'h642e21331397fd28e3911826f15126c62e7c;
       memory[284] = 144'h9c9267c2cedbea090aba5f16f512cdb1a923;
       memory[69] = 144'h7dc504d922f46f27fe6805b1a1ddb4644ad8;
       memory[401] = 144'he3b1026ce10fa54217fd510aa21cfa07edc3;
       memory[564] = 144'h1c496e4e3fb99b2b4fc156df8ab8cd15f6d8;
       memory[466] = 144'h647d696d6c62020a9eb90ae37bee39ba9d1d;
       memory[73] = 144'h5f950e6be2e89b2bf47879b0bf595d52bd26;
       memory[183] = 144'h30a544eb0c7ae907e9a07dbbc389ac2d89d8;
       memory[29] = 144'hfc0502bbb028bf041b606b653f9f125405a8;
       memory[575] = 144'h629944962f263a03ef41c0ddacb6cb4d27e3;
       memory[482] = 144'hf81320a8d086f126e3c2e0bacd78c57afaef;
       memory[489] = 144'h49dc027163ae2e0ed872ae08a448eb7deb34;
       memory[358] = 144'hedea6e9d6eb4f502b5885b9a4c8b0cbf8ede;
       memory[607] = 144'hb0ce49034d174221d889f3ddad83c591342b;
       memory[33] = 144'h51470c731024330f4fb022b36864cde5042d;
       memory[382] = 144'ha94f697c1ee2fa0397c8ba96a5953d72c294;
       memory[107] = 144'h8dfc0222d2e8c6033d226db8140bedaffb90;
       memory[269] = 144'hddcc434d9eb3240c1a4029f939676e8ff71f;
       memory[368] = 144'h3d106606fe65200e2a88672257cc53726a0d;
       memory[58] = 144'hd1c82c8db2950801b71833ef24265717d6ec;
       memory[472] = 144'h77786d864c366d2c4ee1ae6a67480c3f45d1;
       memory[620] = 144'h6ef6650b3d4d270f56591e164eea11e4a086;
       memory[62] = 144'h33d727b9a2872e0f0398772163ee170e934e;
       memory[55] = 144'h906509ee3230d1202fb8db4fd20953ce2dab;
       memory[36] = 144'h15a425c7c0b7d92bc8f0f26bad7107a6299d;
       memory[396] = 144'h975627e9c121412145509e941d40e90be7e3;
       memory[589] = 144'h8b9b481bbdfffa279a59babd92f4462d0d3c;
       memory[574] = 144'h1740635d6f7ef22a0c8146425577747b09d7;
       memory[415] = 144'h8f7308fcb1e0a303969063d2a1be92a8bf27;
       memory[398] = 144'h0fe32f8d8115f723f600bc240e13d568277e;
       memory[494] = 144'hb4d22326b0f7b36fac9da99161322da14417;
       memory[129] = 144'h2d590843715d2423c2da1d460574e9ddb2c7;
       memory[474] = 144'h2dfe684b4c52b222f1d3c6c55d4d3ad0307e;
       memory[478] = 144'he1ac6364ccacf42f4b11c119497e43a2c80d;
       memory[3] = 144'h5dbe0fb390b20901c6506920cbdb5f6e584a;
       memory[61] = 144'hd2f5089a9231472c4ee8a2bc21348f7008f0;
       memory[224] = 144'hef30270370c4ff4dfb852e601b18a67bbdbf;
       memory[180] = 144'h1a0e211cc072c62cd930ba5bfb703e075861;
       memory[46] = 144'h1c3a631afd6b1b02aa0a67380656213c73f1;
       memory[67] = 144'h4aa30a61f27b1123c218ac268f99200b0618;
       memory[570] = 144'hdc4160b72f99b0270dd1ad25bd902661a6ae;
       memory[185] = 144'he8f5489e3ead490e1582d170d43aaa008fb2;
       memory[414] = 144'hdaaa2f5f01934467becd0a699f7fd474aa68;
       memory[556] = 144'h348f6fd56f3e9a26c3d15763fdf7539f9217;
       memory[555] = 144'hfb4d48b73f011c02fb911fec6c00f7ff5822;
       memory[567] = 144'h388248320f536c0ede2167b34d0afbdf5eb2;
       memory[351] = 144'hbfa54c1d0eabdf284bf8c04945711c715f61;
       memory[568] = 144'hc263607e3fc11a2f34f19a646ad3808940eb;
       memory[440] = 144'h35f324ba62528801e5a9cc9614d272e8c225;
       memory[621] = 144'h5ba74e42ddcea12e8f19d24c0d6916cec359;
       memory[236] = 144'hf42622fd42ed0c2f8521a2c4489984daa304;
       memory[232] = 144'hfc3e270ba2dd8b02b56bae7aea553ecb467a;
       memory[218] = 144'h3ea52e6911fcbe4739a5f9973806e688e88b;
       memory[298] = 144'hce816baade9b1a08ad08e6ea81fb6c25d56b;
       memory[176] = 144'h7c292232f0c6082b3fd0c137661be32f44c1;
       memory[27] = 144'h14110832f05047045a303269a590d9fc2dc3;
       memory[481] = 144'h12140c1190ae42058d01262317fbd6a7e779;
       memory[366] = 144'h1ec960c73ec2560a0aa87603b035a91cb921;
       memory[387] = 144'he47542641cf53d63c667f72992a0d3bf38f0;
       memory[251] = 144'he9b10056e0625300a6a3018a2b766083ee65;
       memory[72] = 144'h79ce2a1c72d39808133809ee76c5710e2ce8;
       memory[360] = 144'hf75d66383e2f6f0e0618ad4cf12e6144157a;
       memory[252] = 144'h556024d0d367bb2cdc83c7f861fcb4fd1a6c;
       memory[213] = 144'hd3bd45e09f180f2a461a2abc90fa5e8002c5;
       memory[582] = 144'h19316d84edc5592e0f6386056f4d2bf7cfc9;
       memory[560] = 144'hd7ae69eabf6ba52a8c51af10f45ff1a8ac3d;
       memory[520] = 144'h4bee235ac26d5444eb46a5ada545d3a284aa;
       memory[116] = 144'h2498607b0fe9f449e3259a58c01e216638ec;
       memory[226] = 144'hf5d761a04dabcc485da7939cf2a1d6f46e6f;
       memory[135] = 144'hfd3c0c30c2a3342d096b29fe342ff040a0f3;
       memory[59] = 144'h98a60763f262f2294cc8f22aad2163794354;
       memory[283] = 144'h2e474adceefc3e23c95afe7658a2d7bbbe66;
       memory[240] = 144'h308221a9f28e442ce731f4301ba8b31f617d;
       memory[397] = 144'hde6b0ffb8184ed04bc80a34ade03169ffae8;
       memory[534] = 144'hdddd269ef271e04a8135239c1552432faf75;
       memory[82] = 144'he83f69509f666726c4f235a6c38ac7931297;
       memory[562] = 144'h42bd643c8f2bec24b41143bfece0dc3d10cb;
       memory[289] = 144'h80b54c93ee37382226ca0159c0456cc798c0;
       memory[151] = 144'hd2970203304c7d25af1891a42d9d9844b452;
       memory[331] = 144'h4c3646876ed1a2066812e4c1c2b6d3705259;
       memory[578] = 144'h4d116aad9f434e2fed21799f2600836fa5af;
       memory[416] = 144'hb61165c38c4c4963060d67da8af90091d79d;
       memory[10] = 144'hb01e2dd16090c629c520ef068c95c71f2981;
       memory[91] = 144'h321000038215f6417afc1d3425aa9f9ae315;
       memory[611] = 144'h6b054034cd141c24529997a5601cc2fac642;
       memory[609] = 144'hbb744c97cdd7f82cd91935af8f50bfc596e4;
       memory[171] = 144'h37610e922014750f21400b4da3a7cff3afcb;
       memory[380] = 144'hcde062f16eba320ce2980e80c4cd33f47f60;
       memory[156] = 144'hd6372ff2c0199d230f10c4b991b37428513c;
       memory[206] = 144'hf31165cdbfa28206ecfa9a5f8b11ab8263f4;
       memory[470] = 144'hdbc768552f37ca2b10e3e60b55c3133e4bdb;
       memory[346] = 144'hcafc67425ed768272ef23fc5124d3ea39fbf;
       memory[68] = 144'hdd0623d352dc1c0f8d7885c3d688e7d26ec3;
       memory[355] = 144'hdf7f4c536eac2a207cd853fe7ce3c9ee4834;
       memory[413] = 144'h1a990e185140564b948d37d92bccd9e8cc04;
       memory[405] = 144'h0e970bbed1e6420cd0e0c5758f9acf2ed06f;
       memory[192] = 144'h4cf36b851c249d2f346003d1d030b9cbceb1;
       memory[296] = 144'hada4667bbe8c48096968d0b7aac283c6fe65;
       memory[338] = 144'ha03c6606be6e4a2f2df283d82e523626ed05;
       memory[428] = 144'hbe5d26e24133c1095af930ddd3318a016174;
       memory[529] = 144'h3474075a321c2c6df0d7cafd33dd887d1289;
       memory[467] = 144'h136b4103ac7a6209b9d3c145a0623e7ed2f5;
       memory[204] = 144'h40bd634c5f9cf00e280a3841580061d927d0;
       memory[573] = 144'haf134abebf72390fc2c12abf34a52348a0c0;
       memory[133] = 144'hf20900e441bfa72bac8992f983b809354b47;
       memory[433] = 144'hc55e06d7d3394b2bd7a9bf321f610c20e0fe;
       memory[294] = 144'hab886ec8bc02df09f63a5fca0571296ca45c;
       memory[333] = 144'h63f34b8edeb4380a76f2b4afd531621348bb;
       memory[233] = 144'h3e650229d295990d1391c959e85c010b4b7d;
       memory[8] = 144'hee03232d10be7c21874048e6ed81dc9a4446;
       memory[105] = 144'h78c9443eef24b240ec6f4e76841f3bdc32a5;
       memory[421] = 144'h30e146fd3cecf50f85700c4a56c07cc519e5;
       memory[322] = 144'he00f6300fe5cb123a102c7336437eb530c3d;
       memory[265] = 144'he1cc40e2eec70a0792d0691e5e4a69a40a15;
       memory[14] = 144'hf670207c10562b26d5b0fac3f25d52f4ed09;
       memory[40] = 144'h2a52240920827d08d69a63968ca6d5d5a5c8;
       memory[391] = 144'h3cf508a05144b747502d2be5df81a5b65cd1;
       memory[111] = 144'h47c84cc39f615b0205021a23e902914397c2;
       memory[381] = 144'h9d2545a89e659f2300b836c5d76993a43073;
       memory[164] = 144'h8df227f9d3dff62390e38b97c71debd60a1e;
       memory[616] = 144'hd72063c15d855c0e1369bcfc1dfde29b585c;
       memory[290] = 144'h14e461172ebb7408e8ca6c3f80b64acfdf3b;
       memory[31] = 144'h44b30029906b910c43a0172414a218ab60c2;
       memory[201] = 144'h82a94a593f639f286279b6985614bfefcde2;
       memory[475] = 144'hdede4bf82c71730eb2b393f5957faea1f529;
       memory[56] = 144'hcc0e2d3ce2e2b90a19f88fd4593ce46732ce;
       memory[318] = 144'h0f8665439eeebc261902c5bbf3c235bac787;
       memory[408] = 144'h07d76f278caa6a6b292d828b58acc7df9f66;
       memory[113] = 144'hefb54b540f7c6a0347c2dd5b69eb855e0a35;
       memory[623] = 144'h51fa410d0d5f8300fc9342ad808cd792fcf6;
       memory[63] = 144'h3b160bd2528e91214408403bcab912da0e9b;
       memory[128] = 144'ha470228423adeb02d4ba8cfb10e78c2dfeb5;
       memory[122] = 144'h4ff06bfe9ea0ef4fd99472c47038ae0775f9;
       memory[518] = 144'hcbb963df9cabed4d2484ebb1d5cad3d7938a;
       memory[361] = 144'h896840e1aef79b2f0f384bbd6bab760f0f2b;
       memory[71] = 144'h4be30c96d297ba2c707802ba6cba958f49ec;
       memory[356] = 144'h801c6c5f6e52bb0c717859d6d1f8fe78729f;
       memory[305] = 144'h01734f353e8ccf2da8488a84ad86a9d69066;
       memory[255] = 144'ha14f09a9c3ce1901a89365186fbb6baae2a2;
       memory[324] = 144'h6ee262d0fe135e211772f31ec23804e7e3ee;
       memory[469] = 144'h679047c86fc4560b6f03c354eebb1123033a;
       memory[388] = 144'h3fd9621c5cef8d4f02d7005b7ace9c0fc386;
       memory[379] = 144'h1e3444938ece732546c8db5c248b0d36221f;
       memory[150] = 144'hf56f26f5d0f9ac03ce4852759a2dcd5bb8ca;
       memory[410] = 144'h652a26a281d332271f20d4eab71144fd7488;
       memory[30] = 144'h158f2937301c8e223ee0967fc42b146f2a18;
       memory[158] = 144'hffa32bccd001a9277230ac567cee5e3077c9;
       memory[465] = 144'h093f091ad1fd6b6538c4078cd2f5b8d1da9a;
       memory[327] = 144'hbeaf42e73ea5ca071902602ad726517d210b;
       memory[412] = 144'h5f236d2fec262c6eb6cd281adf28c1ed361e;
       memory[138] = 144'h9672235e31542505f39a1fadef345898677b;
       memory[2] = 144'ha2cd218690c6e72212b0450a82a5281c5229;
       memory[132] = 144'h09022da34148d70ccbc9d7edda0122d53456;
       memory[21] = 144'hb1220dc2e0ccca08b4f0678bd20bdceb9e1e;
       memory[599] = 144'h8ae54ca62d200c28d769731b9abb404fefcf;
       memory[238] = 144'h271d24ee92398f23cea1ba42f02a06cc890a;
       memory[281] = 144'h458a4ae7ce78c52464ba5a25f4b23b5d2ae8;
       memory[300] = 144'hebad6dabfe69970dad78881c70603bbb5c2e;
       memory[9] = 144'h8f300637c07c6b01d7906f5226d43d972142;
       memory[166] = 144'h3dc224cd237fa8297193de4f65076a2e24b8;
       memory[384] = 144'hd9da69a31e06ef0e315840ca95e0e7822b8c;
       memory[155] = 144'h1d1e002c404e1504055379f40ce7c1332020;
       memory[554] = 144'hc5636ee5bfdd392a6091cad1d67e6e10c0b1;
       memory[377] = 144'h5316404fbefbbb27e1a8c2488c5f086d4b99;
       memory[572] = 144'hf4c267b85f1daf2828a16c54d625b1401688;
       memory[191] = 144'had2945204e2222080172c69a2cf1697c68b8;
       memory[604] = 144'h150a6deaddbb620bae8994ceeb6f70a588b6;
       memory[393] = 144'h809b4fa7bc5e3f0043b01c626290239df0a2;
       memory[484] = 144'hdccb2b11b004b02c6732f5f361ae8112aede;
       memory[279] = 144'h117240bf1e8c1d2a12ba13e7593cedb84e5f;
       memory[306] = 144'hfcc26afcde411a0fd1a89f880245e3b391d1;
       memory[513] = 144'hea1445275e4cb82c61a922628f5341920bf8;
       memory[274] = 144'h96fa6fff9e1c5906e3ba178d07fe189d9568;
       memory[553] = 144'h98af4da8bf6f7f0a11e15ea74c6d9e720093;
       memory[595] = 144'haadc497e9d38a22e25998fa36a9de1e89a09;
       memory[121] = 144'h286a40eabd8f5d6d044415606df537c06a53;
       memory[411] = 144'h84780411b156c408fdd084b557bb721e07ca;
       memory[345] = 144'h5d15401cce47b604ede2bec9ea04f78e07da;
       memory[292] = 144'hf8a869de5cf3e800baaa012b25325ec689c6;
       memory[17] = 144'hc9a4014360141b0e404002eb204b1f5dfbd4;
       memory[436] = 144'h41c52a6ac0c4a70c7609daa6dbb3b59b246c;
       memory[275] = 144'h836241256ea96b2b8c9abcb57a224034330e;
       memory[557] = 144'h2d7c483e2f3d000462c1923a156adf41699f;
       memory[458] = 144'hfff029b63198924a54b767dc7328cd15ee8c;
       memory[282] = 144'he97e62812e99c400c37aa492271cb7c00c9d;
       memory[486] = 144'h6f93256fb3581f24f7308928f6ae483bd4b0;
       memory[18] = 144'he68c21b570a3552759c0628e2a96a90dc5fb;
       memory[101] = 144'h13920feab2dd494ae2ff2adee34f5502ff4a;
       memory[225] = 144'ha8af4304adefdf6e65c7bdfe74520a5946c4;
       memory[0] = 144'h43d127a7807e59227cd0c4b49a40917a6c65;
       memory[219] = 144'h48d10b3641bf926f0325f79c48a9b378a1f6;
       memory[342] = 144'h178e6987fe8ca626e912c1218636e37d6e73;
       memory[430] = 144'he71a2653521a4a0ea3ab3f645426ebe47833;
       memory[312] = 144'ha7d168afdee160259492c352e9b79d9f39c1;
       memory[498] = 144'h46b828b433677764acce8c280a4382da6d45;
       memory[449] = 144'h08eb01b7c140666212860abb5fe5ce79e549;
       memory[26] = 144'h1cc120a12030ff263f60d60297feda8bb100;
       memory[90] = 144'h47dd2fedc2d8ab6f946c2f08efc428404bd8;
       memory[487] = 144'h08c402d911d63b03344239d3ce30a1ad454b;
       memory[248] = 144'h550e24549090d3208b7324e7862bd5f34b4a;
       memory[174] = 144'h79362ed7f350412c53f09c19e6c38b32c3f1;
       memory[561] = 144'hfb8240c90f4f470c4361c1c559086bffd782;
       memory[442] = 144'hcc282783c1b3ab0366b9de1ddf2af304277f;
       memory[200] = 144'h12db2631124bb5046ea968bb0d97f8f7d843;
       memory[373] = 144'h04e84ee16e091521bb48c6828964586d2fa5;
       memory[615] = 144'h825c46cbdd436e232bd947832d13f6254b0f;
       memory[367] = 144'h20f74b034e97f1292f480e2ab285d2bbd3d4;
       memory[497] = 144'ha3dc0191838f0f4cef0d0e6b61b9d4de7938;
       memory[521] = 144'h105103e4f28e456ffb66f5a92cfc19a13aca;
       memory[198] = 144'hcb222ee7e01d3d495574e9851c34226b7155;
       memory[325] = 144'h99ab4e9e7e20a3024bc2522dc2be35f6340d;
       memory[93] = 144'h146d44516f18f50b88020d2890333f26398a;
       memory[485] = 144'h773604cc8099880e2c420e8b7a9850ae527c;
       memory[243] = 144'hbeb20c3e92c8940b7f3128a31c57ce2e55d4;
       memory[606] = 144'h29a967c8bdd76708baa9cf744d6a28d4c054;
       memory[610] = 144'h3d7f692abd05810cba59348302c80ad9f462;
       memory[24] = 144'h6b082674801fd02d2630a12d16be27ad9ca8;
       memory[394] = 144'h89d96ae9eca0f66d2b6d954834eb4ab21235;
       memory[451] = 144'h83e30f2d81e6fc654b45bc0f43894394865b;
       memory[261] = 144'hbc314f938e6ca4017ad052e47b1119703e9f;
       memory[343] = 144'hfc3c4e5baec3400b5ac2f16c63eaceb337c7;
       memory[45] = 144'h545a41d67d9dd7282b7a51ff69a67ac4b5bc;
       memory[464] = 144'h37eb20f2c1706e4c55a6d1a64a891246ef6a;
       memory[35] = 144'h42ad0d7d004f99089440ea5d273f77182420;
       memory[499] = 144'h6d10015ac3f7fb4771fe9c94f28785cb95f7;
       memory[54] = 144'hc8f82dcb50bcc102b4aa9b589815d1e1eeb1;
       memory[214] = 144'h5f712b8bf26c15090b797f18a2d1b2beb394;
       memory[266] = 144'ha7886cc20e281b22739006f89a542f1f1241;
       memory[407] = 144'had5a48c4fc00910b55206624c9dbe720f284;
       memory[19] = 144'h8d6c0e4b00e35e0fbd2084c7638a5e9781d7;
       memory[137] = 144'hb36e0fb8a189ac24f4793fb596e2636a26b9;
       memory[100] = 144'hcf1a60f1bf198927118248fbb84aba03522a;
       memory[432] = 144'h05d026f9a023450101fbe62c4a3031b20ba5;
       memory[11] = 144'hdaa90eae40e4a1056f8035ba4b79865fef17;
       memory[558] = 144'h4a3f69d8ff42a725c791152937448e3662dc;
       memory[168] = 144'h62e72bd9c08601267003fad74880a63d11b0;
       memory[519] = 144'h8b8f03f5e1e8da6fe61677517283b129b2e5;
       memory[314] = 144'h9d6164036e26ce2f0632e30573c61d098ee1;
       memory[598] = 144'h4a006f39bdbe950a3d8973fb429adf0a46d0;
       memory[42] = 144'hf64828bef02a8005754a9fbab5e004123ca9;
       memory[612] = 144'h8e7d6440ed29170aa9a9507a592dd9f3c99c;
       memory[476] = 144'h613b652d5ec5db2a2791318581890700637d;
       memory[443] = 144'h4a9e0b9583865d6885e49aeadba25bb19d0b;
       memory[503] = 144'hff630beed0e614424b4ea244b8c667791bbf;
       memory[420] = 144'h3da762a39cffc32a97c0cecb3f91adcde1b6;
       memory[392] = 144'h06cf6cdd5c4b9d2207a0d2ad8557dd95f9a9;
       memory[455] = 144'hc0250a79228ef6636877c735b4abe9ac1b08;
       memory[144] = 144'hb9f4201a3064e80de1090d15c08b01700604;
       memory[592] = 144'h1a58615a3dd42e0b9499bc103adb50b776ef;
       memory[409] = 144'h1d5509a5a1860007b1005d7d8f84952a349a;
       memory[434] = 144'haccc2f6c63bddd05d629e5518df39823731c;
       memory[583] = 144'h44bc444a4d81520274239a80459258a43e82;
       memory[125] = 144'hc16f462d0e6e1d6b9ef7126d6537218c1cd8;
       memory[339] = 144'h12ca4d6f0e2cd6070fc27516e197145da6c7;
       memory[22] = 144'ha51323d5402d422bfb20239bdae68b51f3ca;
       memory[593] = 144'h17bb4edc9de9f4297179fa135c48f675d004;
       memory[178] = 144'he5c92e62b0f6022cb183e5e53e9d2529f592;
       memory[403] = 144'h7f7e4c81dc43cf0ce5900a407c35a0daf836;
       memory[586] = 144'hcbe668a1edba7f006e69b40e10f34b5807da;
       memory[618] = 144'h37e66e429df8ae009ee950047cde44b062a3;
       memory[419] = 144'h6d3e0bfb11559b4cbd2d51d80826f1089fff;
       memory[270] = 144'h3edb6a4a9ea0f02e4130a516e4c06c74ac02;
       memory[471] = 144'h1e094853cfd809061d537f01b9e4c6151776;
       memory[429] = 144'h23660016711fa426e0b92b00516326ade295;
       memory[199] = 144'h5cdc0abb20b0c362b654cfeb9eecd404c6ce;
       memory[532] = 144'hc29862fb7daa0047c026d77067becdff4562;
       memory[76] = 144'hfd452214128d11031bb85337fe8e6a7bf302;
       memory[406] = 144'h860d2db021774a2a064053489dcfa76a04bb;
       memory[165] = 144'hd1d3037c2323a80074138c8cb26ad0816131;
       memory[390] = 144'h711863c09cb7406b9f9d05309f50b165a28c;
       memory[74] = 144'hdec3242a624522029268be6fa10e2172e09f;
       memory[79] = 144'hf1f247354f534e4a3d6fb62c9b6d7a0da696;
       memory[321] = 144'he432444beefc680930220b898b02210479b6;
       memory[181] = 144'h14b2474b6ddf5c0aef42452b0526aa9c7a01;
       memory[264] = 144'hff616388be2b52230920f6f652725bdd3b25;
       memory[431] = 144'h5c3504a5b2dee523005b8c85ad93843ce784;
       memory[566] = 144'hd90f6be59fba13265671eac0dc07de79c85e;
       memory[212] = 144'hbf97661cec7b3c080bc9b5ed270d24a6270f;
       memory[37] = 144'he3f60275809a28044c30a285a7bd2cf6644a;
       memory[509] = 144'h1d250318a32b886034e7e34ec6d913a6fe76;
       memory[126] = 144'h8c0066afee3dfc4c4fb73e4cfc6af41c2ca6;
       memory[145] = 144'h05440417e0c0832f0cea16651cc4e680489d;
       memory[98] = 144'hd2782d35e2676e64ad3f2977f856973ca9fb;
       memory[86] = 144'h07156f748ca9e32ab4f1a9c376f8013ac748;
       memory[246] = 144'hb7492802b21cf624427391dfa2381d46b23b;
       memory[491] = 144'h96d70d1ab3cd5a45e9fd62859227fac7e3b7;
       memory[426] = 144'hc9822a81519c3c2ec7a3d17577dad70875db;
       memory[453] = 144'hc7d30fc671a538609697ffaa63a7f2f8b38d;
       memory[450] = 144'ha3c227d3617c67449345e3e0391962bcb5c0;
       memory[48] = 144'h8a13667c1f10204008e5dc7f82a3ca0efd53;
       memory[38] = 144'h99512ab3506afa08e4fa3603ead6f3e6effd;
       memory[285] = 144'hd9d24405deca3f2eee4aef2322a24025f8ab;
       memory[184] = 144'hdc0561bf4cb46027a25061c492b46e7b8426;
       memory[437] = 144'hc69103c8000552237d69312d5925374496a9;
       memory[328] = 144'h453a6595de08e428ed22737ee93ebbfaad4f;
       memory[417] = 144'h68ce4ed92ca54244791d18f98ef339903e33;
       memory[479] = 144'h79e108ac31cfeb0d6e03e47c2718f9408249;
       memory[490] = 144'h5f8625bef1828a2301c09e35c49045e6ea3a;
       memory[260] = 144'h7c406c58fe08962942b078b00d027f195bff;
       memory[622] = 144'hffa560a2fd750c0268899ede96b16ef41e21;
       memory[15] = 144'hb33c0f12b011010b3b00c1cf26c7f2dadd3e;
       memory[169] = 144'ha4e10ecab0d8d401096356530f8735a55529;
       memory[83] = 144'h42434a5c1c3d1c439fdf901d59f284de6970;
       memory[601] = 144'h13264396cd3d85254eb9a0ccc5f755bac7c6;
       memory[585] = 144'h04b54b321d1bd8228b79df9b0731b47156bc;
       memory[454] = 144'h70202a05a25a0144d8752ef2d3adb5193917;
       memory[262] = 144'h623266a75e26be23ed6047e644c1f93d3405;
       memory[263] = 144'h8fe641d11ec5a105f3d0ad75319ad68e11c5;
       memory[386] = 144'h0a6367c94e949b0ed78a782688f6aaf2bb2b;
       memory[383] = 144'he30141d26eaa622b7508cf5d3ddb085e4f2d;
       memory[25] = 144'hdb860bccf02e5b09c7f0bf4f32194b94f2df;
       memory[579] = 144'h25fa4853ffcf3b01e8e1de410e639a4ebcbd;
       memory[541] = 144'h72f44aa0ff24d52ca21864149d2f780046dc;
       memory[577] = 144'hc5c94e28cfc75f000981ee9a3228e81eded4;
       memory[603] = 144'hbe774c92ada1212a7fc98013e3e0ff0dd57d;
       memory[12] = 144'hfb4f2c783024eb2cb630a10b08bb801c8f1a;
       memory[348] = 144'h85aa68212e7ce9290f22a493a96542404fe5;
       memory[202] = 144'h696b62380ff2f908d2f998c0352dc5d80db8;
       memory[344] = 144'h32786ebecefb4724b042dfd115b6e9f4715b;
       memory[522] = 144'h4c7d25eb11f54f4458264911d5a90013fb20;
       memory[197] = 144'h2cf206ece0ac4c66f0c407444ce8c8c02f0a;
       memory[444] = 144'ha39d236ad3e104091b39b3437a1676a9df0d;
       memory[182] = 144'h48b7694a7f39e426f59097c0397e862bf90d;
       memory[504] = 144'hb868207710c0036ae3fd2fda422d4942549d;
       memory[337] = 144'h979741189ee89d09ebf2887f857f711600f5;
       memory[329] = 144'h2389402cde93390ea5b207c12bec1544d0dc;
       memory[316] = 144'h204068248e04802481e26a10260652574a40;
       memory[1] = 144'hdb620da0d052e80e06c0534e5f328e7f3c25;
       memory[614] = 144'he8cc64d82d41b703dc7952a5efa65062dac2;
       memory[334] = 144'ha56e6226beda312127d21091beecbeaf8f39;
       memory[374] = 144'hdd2f6edf3ef25f06df283d6ada1031adabac;
       memory[495] = 144'h71820d24738fb843801d073ddbb957f5b45b;
       memory[395] = 144'hed4501b571ba93076f90f9ffa1e0d7d9fab1;
       memory[210] = 144'h5b15618ddc81ef06d3e99d6dc439f906b969;
       memory[41] = 144'h92560b5f4091ef2db2eac652b6f50328c57c;
       memory[222] = 144'h279a6a5b6d94b107dc8a8e10ade86e2ee9db;
       memory[286] = 144'h1c0e6fcfbea6ec01826a00e06c67d5772bd5;
       memory[594] = 144'h003460750d23e40d7a791648d67e2ccba843;
       memory[23] = 144'hec900dc200304f06cb90b7b8c6914e26803c;
       memory[16] = 144'h3a7424faf0c0b2222790918ae23d50c2e491;
       memory[493] = 144'hd13408c0c0996942cefd2a2e03fab2d6d847;
       memory[552] = 144'hc81363558fdebe2f7f715aafc22d19cc68cc;
       memory[350] = 144'h95516d211ec4c40bc5789961d0dbefdcdfee;
       memory[515] = 144'h3d994f663e8a462744f99f56ad139f87d875;
       memory[547] = 144'hd3a243248fa8930d79c1366250593bf7bd96;
       memory[613] = 144'h24884877cd11b122f709bc7c3ca346cb3c03;
       memory[134] = 144'h5ba424cf7102a700cdf916766fd205f82ba0;
       memory[277] = 144'h312742027ecbe521c41a0dd97375acd27284;
       memory[267] = 144'h65cc407e0e04b40fae2035e0ead50440ea13;
       memory[84] = 144'h4286261441f66c6d549f5304d18648e15eb7;
       memory[5] = 144'h7fbe0bea503c580032a0e15a3cafeda921a9;
       memory[531] = 144'hb2da42ce9faa636a0815d24394c2fbdb7b1e;
       memory[591] = 144'hc37142be4dc1bb242e798d198e10639e9620;
       memory[280] = 144'hbdde6194aeef4c0be66a8dbb678535d5288b;
       memory[539] = 144'hc1c20fc74022286e3705397ddee2fcb69607;
       memory[189] = 144'h6ca047b4ae4ad646ea1f8e1e0ec9e23006c1;
       memory[605] = 144'h2c7c494c3d55bb29d269ab4a8ffb23b781ab;
       memory[75] = 144'h941804ac52987b2bd638263b3ab96d0a7681;
       memory[205] = 144'h5cff4a6c7fa7332a40da06434c271664591f;
       memory[543] = 144'h12cb4d510f9cbe2b57cb12d6b6a441dc044c;
       memory[159] = 144'h00830f0380551204c430ee7bb4edf296a8a1;
       memory[60] = 144'h40f529f7524f4605079892fb197eedace033;
       memory[190] = 144'h0e3e6a718ebe946f88af3dd633b056c56b58;
       memory[551] = 144'h9c654f102f858f05b43197558b5582e85e61;
       memory[148] = 144'hfdf7270d1058060a9228a7945bb39d1aa726;
       memory[362] = 144'hd51d641c8e609c0bc17898a98786c75e3528;
       memory[142] = 144'hbba12aafa3ae41062819796c6fa09a88cd29;
       memory[81] = 144'h0bec0e3f82499146664f7d05f31dadcbda8f;
       memory[315] = 144'ha6634b404ef3940341329110340b9978eeea;
       memory[528] = 144'h3d0a67996f4a3008eeaa68e30aedea14f240;
       memory[288] = 144'ha85c69df0edffd03b24aca7e1d837a76cfe9;
       memory[44] = 144'h0ba062d9bdb6c60c6deab3429cd605f17b02;
       memory[106] = 144'h6fc26768ff9a2966d77fccc39d169596a200;
       memory[559] = 144'he4f94e376fb45b0f8b6115469e2f9bde0c89;
       memory[456] = 144'h862c292551c13b4708e7b0e22cec5ac0b3ff;
       memory[550] = 144'h71a16352bfa6f8260321738778fe6b961d64;
       memory[511] = 144'h497b08800128d265c2b4d707344695df0a23;
       memory[64] = 144'hbf8820a6e2700c05999806b6ac4ad4c7226b;
       memory[571] = 144'haa2448b04ff3a50b7801a827a6b1523934ff;
       memory[85] = 144'hfec600bf4141a70986525ce40e6868041884;
       memory[250] = 144'h8d092e4f2030122a89334364c6eb52be25fb;
       memory[452] = 144'hf8012417117d6848f4f7803c3d539182d8b5;
       memory[548] = 144'h959267681f85b22372e100344b8123c40f6d;
       memory[124] = 144'hf69a63617ed75f4291a454025673db15d55b;
       memory[597] = 144'h7be84f940d31532c10c94e40774fddd53d5b;
       memory[590] = 144'h7ebe6d16bda39900a639231d85a373629519;
       memory[524] = 144'h0dbc26a6c22f1f458416da6a5aee6bde732b;
       memory[20] = 144'h535f299540f73a2b5d90548873d9fd9f7a56;
       memory[53] = 144'h5adf0c3a007e6b6b9ac78310e6ecbbae08f7;
       memory[372] = 144'hb33f613f2e401e0641b8778fc93eb52e59cd;
       memory[227] = 144'h96054e62cdc1386c02a76a6697cb67454e56;
       memory[371] = 144'hf6d743c35e4aae248ff8c5ec6b081bb17304;
       memory[6] = 144'h2e35225810e72f28d440763ce7258725d280;
       memory[544] = 144'hf37a6935df60ee09760bbbd4ef1958c46b18;
       memory[445] = 144'h2e0f0c4b2325216935542798a5f0e8f169a9;
       memory[308] = 144'h4aeb69495ec89a09f5f8e480d4ccc2e82e9f;
       memory[50] = 144'h78656b526f7a7e41a17516d0e01c2048eef3;
       memory[459] = 144'h989c040c71da1d60c7f426ce9ab729454090;
       memory[457] = 144'hec1509d981dd7863f3049a6a9f0b2800bb64;
       memory[538] = 144'h657823bf9262834907e6cc928f458392b6ab;
       memory[512] = 144'h01d167ba5c9e6a0d6b294b238cfa402d24e2;
       memory[584] = 144'hfc5e6d8dad16b00c70299531ebdedf42d1ad;
       memory[78] = 144'hee942555c2de6f2ac35263c8272686749f01;
       memory[507] = 144'h497f002f40df996c1b57370825ec7b3c7ad0;
       memory[301] = 144'hd06e4075ce618d2eab18f8e742b76901591c;
       memory[354] = 144'h90346fddaec2ec0090482cf0f1746abf95b8;
       memory[157] = 144'h17480aa750743c02c2e02f70aa5c8c7cd7a1;
       memory[477] = 144'h24f743945c4f9b0d6dd18681fa2eb338b541;
       memory[245] = 144'h08ce0b7ed2ef0809c16195c6cdb3dc69b4d0;
       memory[527] = 144'h448a46a63f027a27c3d819cac8c6d1053996;
       memory[149] = 144'h86f706c5f0bc6d2c6bf8ad0cebe353e0e650;
       memory[57] = 144'h0cae0c4ba2deab2911480b3e48f979449e77;
       memory[506] = 144'h43b9249d0034e140dcc7e41d8ef5da813572;
       memory[488] = 144'h058e27c133a3f225dcc22b98b085d6b8d15c;
       memory[242] = 144'h0d3f20b372dccc23413195450db112e1d7b2;
       memory[502] = 144'he89e221c70072164748e169c549765277d36;
       memory[244] = 144'ha13d29eaf226d32bca6161641eb84b47207c;
       memory[546] = 144'h85a16b14afcde3216121a94af62cbccd54f4;
       memory[463] = 144'h816302e2e1e71a611236ac30fd84464e595d;
       memory[65] = 144'h90850c87827ecb22e2a836a41a8a8d18b864;
       memory[130] = 144'h2a8e2f89e1bdce0ba06a0af1c864fff9b3ba;
       memory[602] = 144'h65c16da7dddf4c0183e9d5fd8455bf4cff7e;
       memory[154] = 144'h2a362670f04e260abf695d6755c2c5d05f0f;
       memory[237] = 144'h41600564c2f6a0044d51e31699b5cafeb899;
       memory[619] = 144'h61e2451f0d690d23c9e96c0294b9ac85b67b;
       memory[80] = 144'hf29b273e327e786cad4f19479b1f6f67fd9d;
       memory[357] = 144'h03794f1b5e5fc520e4b82be6143a849942ef;
       memory[535] = 144'hff21064bd2c006619b360aa2a3e08e8aca1a;
       memory[299] = 144'hd8dd481ebe782c2ca9980aa66f2119c28a5b;
       memory[364] = 144'he4026f92aeaeb301c8481917dfd2ce137f82;
       memory[47] = 144'h6f4f427b0dac9667d0779520ae9660bf5722;
       memory[253] = 144'h92430236c3c4e703ec13a214d3590e487d14;
       memory[160] = 144'h2b302c8780958f2aceb02567ddd0a5ac42c3;
       memory[462] = 144'h3e50220a623ddc4ba416929872540132f9e6;
       memory[51] = 144'h0dde07706217516416f7363c58f1c2f77448;
       memory[118] = 144'h8d4561980dc88842c89615c2f47b9d7c0da1;
       memory[216] = 144'hafd126b7f0cccd05407b1da8984779ef4fdc;
       memory[370] = 144'hfb886127aefd4409b1987ba09f05596396f6;
       memory[92] = 144'h8ff92008c2d8b42a9dd1a2b42a2be2a718b8;
       memory[39] = 144'h64550cc7e0bc9726576a043c1b44e8329e65;
       memory[258] = 144'h86fa6b3bbe5a6b20663061c6cd4a3a0ac7fa;
       memory[152] = 144'h57382c34e08dc50aa31ac76d7d15b0296d39;
       memory[302] = 144'h027565178eb6ed06cb08d5f4333b978b55ab;
       memory[293] = 144'h128e48c13c0b782e345a4e1cd9b59e45b5de;
       memory[141] = 144'hc9d40a8951dc222734e9dac6e9e40ff12145;
       memory[268] = 144'h900d6800dedb4421e120649e94f88a13111d;
       memory[441] = 144'h45dd031da2431222cf49a684430f34104050;
       memory[211] = 144'h8e0d4e073c486a2e12c9daf54b57fb43182b;
       memory[103] = 144'hf93b0f487281080446b27e112576344700b2;
       memory[231] = 144'h0262018c70a59520005854efeed3a98dd955;
       memory[525] = 144'h83780e27a0a6086cfc45d928c1bc017ba567;
       memory[115] = 144'h8d4c40f91fa98a4ab0cf85431795fda8109d;
       memory[207] = 144'he58547baac0209246cca0e9aa6da3e7642df;
       memory[596] = 144'h6d666e55bd81ba0e34e9689143151d837dde;
       memory[399] = 144'hf41d0922d1b50d029520e4ff4a5755d63ba6;
       memory[517] = 144'hf66a419bee28ad241a6986d2fabda7f65815;
       memory[127] = 144'h8b9643d04ef51b6d20d72b8ef5a02963e8b6;
       memory[175] = 144'h1816042ce37cb5031e908416fd5c51f77c0c;
       memory[119] = 144'ha2fc4df6bd9b516175344c7e89b702deecb1;
       memory[195] = 144'hadf445a31eea15235cfb000c9c7043b29633;
       memory[278] = 144'h71676afd2e9e3f04efbae808530ec42f3e9a;
       memory[422] = 144'hd536602b1c898a63543d6c0d6acd663c5e3b;
       memory[447] = 144'h7ce30caa6259f662e4762f038ce657fddabc;
       memory[87] = 144'h16170cf601289244fe3c879a5be1fc84b7d1;
       memory[365] = 144'had854ba4be80332c4a28b0009e7f83a88585;
       memory[203] = 144'hc3704372df59ac20e7cacc26df9781fd24ef;
       memory[533] = 144'head20a8a70f30968d4458a20f290e2f91362;
       memory[438] = 144'ha07b21a8c0c8a9074dd936c157eceb340e4d;
       memory[170] = 144'h3901271730b93322a2938b0d1406bcf2b4a3;
       memory[109] = 144'h226a46983fe5a805869214420706a3fe9b4d;
       memory[173] = 144'h541b05920016230486803d6e79787af45bac;
       memory[569] = 144'h6e7a42b51f807e01d3410aa16a461bc7fdef;
       memory[435] = 144'h0f9606b470d90b2012195271df4fe7efdb4b;
       memory[4] = 144'h54902f3040b4cc2991d0766847dc02547898;
       memory[235] = 144'haa40059ce2d8560a7811468d3e1872484cb9;
       memory[140] = 144'hd81526a71143d9096619067f41f3b1a7104f;
       memory[508] = 144'hf91b276af3bc0742a7d742fb0d45c86a786b;
       memory[461] = 144'h0d0f0e1df22fb961e7166a0aa826d8d28ce1;
       memory[423] = 144'ha1040732d1d53400e9b0755d1c05507eb769;
       memory[500] = 144'hc0702989e0d25d6765fc4fbbb014238c79ea;
       memory[186] = 144'h944b6b237c2e3263e67f45eb7a27455f3087;
       memory[94] = 144'hf2a524ee723dbe6fdfafa127c4ceaac9301d;
       memory[97] = 144'hfb2303f472e3c949a60fca2bda96ce59475f;
       memory[163] = 144'hcd8f0c2f03c2af0eb880888124435b2729cf;
       memory[310] = 144'haa366f0d0e1a1809f4d8f19c736a343c60d7;
       memory[501] = 144'h007b0c0eb245b34bd80e5bf0f1d13501612d;
       memory[153] = 144'h4f110ac7c07f3e2f538a2181008bf388a238;
       memory[496] = 144'hb2d02ea193f3ae6c88deab740f5b0d40abe6;
       memory[330] = 144'hed306ac13e3b0a23b1627839028642a6f0a2;
       memory[104] = 144'h6315626fcfbf5962fd2fd6516cbbf2198cfa;
       memory[341] = 144'hd96a442bbe672c0d210206ca745589f6e521;
       memory[221] = 144'h48b24bf9fe4ced23a6ba3ba78bb9b1eace0b;
       memory[220] = 144'hc88e2e9083d9dc061688095b73a1989ec0f6;
       memory[309] = 144'h2d3047f6ae5fa02d5ee8a06907667b3874d0;
       memory[271] = 144'h0a884679ae1d3e048ee0247efc0271912c85;
       memory[404] = 144'hb41820cc81f7da2e06802dd29cf58174a5d6;
       memory[161] = 144'h07c104120313090c087057b3a6ac31439d45;
       memory[223] = 144'hc17b4da95d50462b1ac8776c781f57a8e41c;
       memory[587] = 144'hcdef4cb78dca002521e9b21013bd70b6b3a0;
       memory[234] = 144'h51812459624f7222fae111da0d0850bdebba;
       memory[13] = 144'h00760944b015fc0f9f70cb28dddcb1472016;
       accumulator = 0;
   end
   
   reg [15:0] accumulator;
   always @(posedge clk) begin
       graphicsMem[counter] = accumulator^result[counter];
       accumulator = result[counter];
       counter = #1 counter + 1;
   end
endmodule

module generator(in, count, counter, out, vb);
   input [143:0] in;
   input [31:0]  counter, count;
   output [15:0] out;
   output 	 vb;
   reg 		 outMem;
   wire 	 outMemInternal;
   
   initial outMem = 0;
   assign outMemInternal = count == counter ? 1'b1 : 1'b0;
   always @(outMemInternal) outMem = ~outMem;
   assign vb = ~outMem;
   assign out = (count == counter) ? {{in[127:124]},{in[107:104]},{in[87:84]},{in[67:64]}} : {{2{in[44-:2]}},{2{in[40-:2]}},{2{in[36-:2]}},{2{in[32-:2]}}};
endmodule
